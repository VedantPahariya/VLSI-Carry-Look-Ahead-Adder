magic
tech scmos
timestamp 1731482030
<< nwell >>
rect -261 314 -229 351
rect -202 314 -177 330
rect -261 310 -177 314
rect -261 295 -178 310
rect -261 259 -202 295
rect -217 256 -202 259
rect -165 226 -145 267
rect -210 143 -178 180
rect 16 173 28 176
rect -210 88 -151 143
rect 4 141 28 173
rect -129 96 -94 120
rect 44 105 64 146
rect -166 85 -151 88
rect -114 55 -94 96
<< ntransistor >>
rect -191 279 -189 289
rect -250 213 -248 253
rect -242 213 -240 253
rect -175 254 -171 256
rect -223 210 -221 250
rect -215 210 -213 250
rect -175 238 -171 240
rect 15 125 17 135
rect 34 133 38 135
rect 34 117 38 119
rect -145 107 -135 109
rect -199 42 -197 82
rect -191 42 -189 82
rect -124 83 -120 85
rect -172 39 -170 79
rect -164 39 -162 79
rect -124 67 -120 69
<< ptransistor >>
rect -250 265 -248 345
rect -242 265 -240 345
rect -223 268 -221 308
rect -215 268 -213 308
rect -191 301 -189 321
rect -159 254 -151 256
rect -159 238 -151 240
rect -199 94 -197 174
rect -191 94 -189 174
rect 15 147 17 167
rect -172 97 -170 137
rect -164 97 -162 137
rect 50 133 58 135
rect 50 117 58 119
rect -123 107 -103 109
rect -108 83 -100 85
rect -108 67 -100 69
<< ndiffusion >>
rect -196 283 -191 289
rect -192 279 -191 283
rect -189 285 -188 289
rect -189 279 -184 285
rect -251 249 -250 253
rect -255 213 -250 249
rect -248 217 -242 253
rect -248 213 -247 217
rect -243 213 -242 217
rect -240 249 -239 253
rect -175 256 -171 257
rect -175 253 -171 254
rect -240 213 -235 249
rect -228 214 -223 250
rect -224 210 -223 214
rect -221 210 -215 250
rect -213 246 -212 250
rect -213 210 -208 246
rect -175 240 -171 241
rect -175 237 -171 238
rect 34 135 38 136
rect 10 129 15 135
rect 14 125 15 129
rect 17 131 18 135
rect 17 125 22 131
rect 34 132 38 133
rect 34 119 38 120
rect 34 116 38 117
rect -141 110 -135 114
rect -145 109 -135 110
rect -145 106 -135 107
rect -145 102 -139 106
rect -200 78 -199 82
rect -204 42 -199 78
rect -197 46 -191 82
rect -197 42 -196 46
rect -192 42 -191 46
rect -189 78 -188 82
rect -124 85 -120 86
rect -124 82 -120 83
rect -189 42 -184 78
rect -177 43 -172 79
rect -173 39 -172 43
rect -170 39 -164 79
rect -162 75 -161 79
rect -162 39 -157 75
rect -124 69 -120 70
rect -124 66 -120 67
<< pdiffusion >>
rect -255 269 -250 345
rect -251 265 -250 269
rect -248 265 -242 345
rect -240 341 -239 345
rect -240 265 -235 341
rect -192 317 -191 321
rect -224 304 -223 308
rect -228 268 -223 304
rect -221 272 -215 308
rect -221 268 -220 272
rect -216 268 -215 272
rect -213 304 -212 308
rect -213 268 -208 304
rect -196 301 -191 317
rect -189 305 -184 321
rect -189 301 -188 305
rect -155 257 -151 261
rect -159 256 -151 257
rect -159 253 -151 254
rect -155 249 -151 253
rect -155 241 -151 245
rect -159 240 -151 241
rect -159 237 -151 238
rect -154 233 -151 237
rect -204 98 -199 174
rect -200 94 -199 98
rect -197 94 -191 174
rect -189 170 -188 174
rect -189 94 -184 170
rect 14 163 15 167
rect 10 147 15 163
rect 17 151 22 167
rect 17 147 18 151
rect -173 133 -172 137
rect -177 97 -172 133
rect -170 101 -164 137
rect -170 97 -169 101
rect -165 97 -164 101
rect -162 133 -161 137
rect -162 97 -157 133
rect 54 136 58 140
rect 50 135 58 136
rect 50 132 58 133
rect 54 128 58 132
rect 54 120 58 124
rect 50 119 58 120
rect -123 110 -107 114
rect 50 116 58 117
rect 55 112 58 116
rect -123 109 -103 110
rect -123 106 -103 107
rect -119 102 -103 106
rect -104 86 -100 90
rect -108 85 -100 86
rect -108 82 -100 83
rect -104 78 -100 82
rect -104 70 -100 74
rect -108 69 -100 70
rect -108 66 -100 67
rect -103 62 -100 66
<< ndcontact >>
rect -196 279 -192 283
rect -188 285 -184 289
rect -255 249 -251 253
rect -247 213 -243 217
rect -239 249 -235 253
rect -175 257 -171 261
rect -228 210 -224 214
rect -212 246 -208 250
rect -175 249 -171 253
rect -175 241 -171 245
rect 34 136 38 140
rect 10 125 14 129
rect 18 131 22 135
rect 34 128 38 132
rect 34 120 38 124
rect -145 110 -141 114
rect -139 102 -135 106
rect -204 78 -200 82
rect -196 42 -192 46
rect -188 78 -184 82
rect -124 86 -120 90
rect -177 39 -173 43
rect -161 75 -157 79
rect -124 78 -120 82
rect -124 70 -120 74
<< pdcontact >>
rect -255 265 -251 269
rect -239 341 -235 345
rect -196 317 -192 321
rect -228 304 -224 308
rect -220 268 -216 272
rect -212 304 -208 308
rect -188 301 -184 305
rect -159 257 -155 261
rect -159 249 -155 253
rect -159 241 -155 245
rect -204 94 -200 98
rect -188 170 -184 174
rect 10 163 14 167
rect 18 147 22 151
rect -177 133 -173 137
rect -169 97 -165 101
rect -161 133 -157 137
rect 50 136 54 140
rect 50 128 54 132
rect 50 120 54 124
rect -107 110 -103 114
rect -123 102 -119 106
rect -108 86 -104 90
rect -108 78 -104 82
rect -108 70 -104 74
<< polysilicon >>
rect -250 345 -248 348
rect -242 345 -240 348
rect -191 321 -189 324
rect -223 308 -221 311
rect -215 308 -213 311
rect -191 289 -189 301
rect -191 276 -189 279
rect -250 261 -248 265
rect -250 253 -248 256
rect -242 253 -240 265
rect -223 250 -221 268
rect -215 260 -213 268
rect -215 250 -213 255
rect -178 254 -175 256
rect -171 255 -168 256
rect -163 255 -159 256
rect -171 254 -159 255
rect -151 254 -148 256
rect -250 210 -248 213
rect -242 210 -240 213
rect -179 238 -175 240
rect -171 238 -168 240
rect -162 238 -159 240
rect -151 238 -150 240
rect -223 207 -221 210
rect -215 207 -213 210
rect -199 174 -197 177
rect -191 174 -189 177
rect 15 167 17 170
rect -172 137 -170 140
rect -164 137 -162 140
rect 15 135 17 147
rect 31 133 34 135
rect 38 134 41 135
rect 46 134 50 135
rect 38 133 50 134
rect 58 133 61 135
rect 15 122 17 125
rect 29 117 34 119
rect 38 117 41 119
rect 47 117 50 119
rect 58 117 59 119
rect -148 107 -145 109
rect -135 107 -123 109
rect -103 107 -100 109
rect -199 90 -197 94
rect -199 82 -197 85
rect -191 82 -189 94
rect -172 79 -170 97
rect -164 89 -162 97
rect -164 79 -162 84
rect -127 83 -124 85
rect -120 84 -117 85
rect -112 84 -108 85
rect -120 83 -108 84
rect -100 83 -97 85
rect -199 39 -197 42
rect -191 39 -189 42
rect -128 67 -124 69
rect -120 67 -117 69
rect -111 67 -108 69
rect -100 67 -99 69
rect -172 36 -170 39
rect -164 36 -162 39
<< polycontact >>
rect -195 290 -191 294
rect -240 260 -236 264
rect -227 260 -223 264
rect -183 238 -179 242
rect -150 238 -146 242
rect 11 136 15 140
rect 25 117 29 121
rect 59 117 63 121
rect -134 109 -130 113
rect -189 89 -185 93
rect -176 89 -172 93
rect -132 67 -128 71
rect -99 67 -95 71
<< metal1 >>
rect -261 349 -228 352
rect -238 345 -235 349
rect -231 305 -228 349
rect -212 327 -177 330
rect -212 308 -208 327
rect -196 321 -193 327
rect -224 305 -212 308
rect -201 311 -160 314
rect -201 294 -198 311
rect -187 296 -184 301
rect -201 291 -195 294
rect -235 288 -198 291
rect -187 293 -177 296
rect -187 289 -184 293
rect -259 265 -255 268
rect -259 253 -256 265
rect -235 264 -232 288
rect -196 276 -193 279
rect -202 273 -188 276
rect -219 266 -216 268
rect -236 261 -227 264
rect -219 263 -205 266
rect -259 250 -255 253
rect -251 250 -239 253
rect -208 247 -205 263
rect -211 239 -208 246
rect -260 236 -208 239
rect -247 209 -244 213
rect -228 209 -224 210
rect -202 209 -199 273
rect -181 267 -177 293
rect -182 264 -177 267
rect -164 266 -160 311
rect -182 261 -179 264
rect -164 263 -147 266
rect -159 261 -155 263
rect -182 258 -175 261
rect -182 242 -179 258
rect -171 249 -159 252
rect -169 245 -166 249
rect -171 242 -159 245
rect -167 228 -164 242
rect -150 242 -147 263
rect -256 206 -199 209
rect -210 178 -177 181
rect -187 174 -184 178
rect -180 134 -177 178
rect 4 173 28 176
rect 10 167 13 173
rect 5 157 54 160
rect 5 140 8 157
rect 19 142 22 147
rect 51 145 54 157
rect 51 142 62 145
rect 19 140 29 142
rect 51 140 54 142
rect 5 137 11 140
rect -173 134 -161 137
rect -157 134 -151 137
rect 19 139 34 140
rect 19 135 22 139
rect -154 126 -151 134
rect 26 137 34 139
rect -154 123 -104 126
rect -184 119 -130 120
rect -184 117 -110 119
rect -208 94 -204 97
rect -208 82 -205 94
rect -184 93 -181 117
rect -133 116 -110 117
rect -151 111 -145 114
rect -168 95 -165 97
rect -185 90 -176 93
rect -168 92 -154 95
rect -208 79 -204 82
rect -200 79 -188 82
rect -157 76 -154 92
rect -160 68 -157 75
rect -207 65 -157 68
rect -196 38 -193 42
rect -177 38 -173 39
rect -151 38 -148 111
rect -133 113 -130 116
rect -135 102 -123 105
rect -131 90 -128 102
rect -113 95 -110 116
rect -107 114 -104 123
rect 10 122 13 125
rect 10 119 22 122
rect 26 121 29 137
rect 38 128 50 131
rect 40 124 43 128
rect 38 121 50 124
rect 42 107 45 121
rect 59 121 62 142
rect -113 92 -96 95
rect -108 90 -104 92
rect -131 87 -124 90
rect -131 71 -128 87
rect -120 78 -108 81
rect -118 74 -115 78
rect -120 71 -108 74
rect -116 57 -113 71
rect -99 71 -96 92
rect -205 35 -148 38
<< pm12contact >>
rect -253 256 -248 261
rect -217 255 -212 260
rect -168 255 -163 260
rect -202 85 -197 90
rect -166 84 -161 89
rect 41 134 46 139
rect -117 84 -112 89
<< pdm12contact >>
rect -159 232 -154 237
rect 50 111 55 116
rect -108 61 -103 66
<< ndm12contact >>
rect -176 232 -171 237
rect 33 111 38 116
rect -125 61 -120 66
<< metal2 >>
rect -248 256 -217 259
rect -212 256 -168 259
rect -166 236 -163 255
rect -171 233 -159 236
rect 2 153 44 156
rect 41 139 44 153
rect 43 115 46 134
rect 38 112 50 115
rect -197 85 -166 88
rect -161 85 -117 88
rect -115 65 -112 84
rect -120 62 -108 65
use XOR  XOR_0
timestamp 1731446490
transform 1 0 274 0 1 237
box -351 -83 -274 -26
<< labels >>
rlabel metal1 -188 36 -188 36 1 gnd
rlabel metal1 -190 180 -190 180 5 VDD
rlabel metal1 -206 86 -206 86 3 out
rlabel metal1 -182 91 -182 91 7 A
rlabel metal2 -182 86 -182 86 7 B
rlabel metal1 43 108 43 108 3 out
rlabel metal1 12 175 12 175 5 VDD
rlabel metal1 15 120 15 120 1 gnd
rlabel metal1 7 138 7 138 1 A
rlabel metal1 -115 58 -115 58 3 out
rlabel metal1 -132 117 -132 117 3 A
rlabel metal1 -150 109 -150 109 3 gnd
rlabel metal1 -166 229 -166 229 3 out
rlabel metal2 -233 257 -233 257 7 B
rlabel metal1 -233 262 -233 262 7 A
rlabel metal1 -257 257 -257 257 3 out
rlabel metal1 -241 351 -241 351 5 VDD
rlabel metal1 -239 207 -239 207 1 gnd
rlabel metal1 -199 292 -199 292 1 A
rlabel metal1 -191 274 -191 274 1 gnd
rlabel metal1 -194 329 -194 329 5 VDD
<< end >>
