magic
tech scmos
timestamp 1731409263
<< nwell >>
rect -82 43 -30 69
rect -82 17 19 43
rect -30 11 19 17
<< ntransistor >>
rect -18 49 -16 69
rect -12 49 -10 69
rect 6 49 8 69
rect 12 49 14 69
rect -71 0 -69 11
rect -49 0 -47 11
<< ptransistor >>
rect -71 23 -69 63
rect -65 23 -63 63
rect -49 23 -47 63
rect -43 23 -41 63
rect -18 17 -16 37
rect 6 17 8 37
<< ndiffusion >>
rect -24 56 -18 69
rect -19 51 -18 56
rect -24 49 -18 51
rect -16 49 -12 69
rect -10 53 -4 69
rect -10 49 -8 53
rect 0 56 6 69
rect 5 51 6 56
rect 0 49 6 51
rect 8 49 12 69
rect 14 53 20 69
rect 14 49 16 53
rect -76 4 -71 11
rect -72 0 -71 4
rect -69 7 -68 11
rect -69 0 -64 7
rect -54 4 -49 11
rect -50 0 -49 4
rect -47 7 -46 11
rect -47 0 -42 7
<< pdiffusion >>
rect -72 59 -71 63
rect -76 23 -71 59
rect -69 23 -65 63
rect -63 27 -58 63
rect -63 23 -62 27
rect -50 59 -49 63
rect -54 23 -49 59
rect -47 23 -43 63
rect -41 27 -36 63
rect -41 23 -40 27
rect -23 23 -18 37
rect -19 19 -18 23
rect -23 17 -18 19
rect -16 33 -15 37
rect -16 17 -11 33
rect 1 23 6 37
rect 5 19 6 23
rect 1 17 6 19
rect 8 33 9 37
rect 8 17 13 33
<< ndcontact >>
rect -8 49 -4 53
rect 16 49 20 53
rect -76 0 -72 4
rect -68 7 -64 11
rect -54 0 -50 4
rect -46 7 -42 11
<< pdcontact >>
rect -76 59 -72 63
rect -62 23 -58 27
rect -54 59 -50 63
rect -40 23 -36 27
rect -23 19 -19 23
rect -15 33 -11 37
rect 1 19 5 23
rect 9 33 13 37
<< polysilicon >>
rect -71 63 -69 66
rect -65 63 -63 74
rect -49 63 -47 66
rect -43 63 -41 70
rect -18 69 -16 73
rect -12 69 -10 70
rect 6 69 8 73
rect 12 69 14 70
rect -18 37 -16 49
rect -12 46 -10 49
rect 6 37 8 49
rect 12 46 14 49
rect -71 11 -69 23
rect -65 20 -63 23
rect -49 11 -47 23
rect -43 20 -41 23
rect -18 14 -16 17
rect 6 14 8 17
rect -71 -3 -69 0
rect -49 -3 -47 0
<< polycontact >>
rect -63 70 -59 74
rect -44 70 -40 74
rect -12 70 -8 74
rect 12 70 16 74
rect 2 44 6 48
rect -75 12 -71 16
rect -53 12 -49 16
rect -22 12 -18 16
<< metal1 >>
rect -59 71 -44 74
rect -40 71 -12 74
rect -8 71 12 74
rect -75 64 -27 67
rect -75 63 -72 64
rect -54 63 -50 64
rect -61 16 -58 23
rect -39 16 -36 23
rect -30 23 -27 64
rect -7 47 -4 49
rect -7 44 2 47
rect 17 47 20 49
rect 17 44 26 47
rect -7 37 -4 44
rect 17 37 20 44
rect -11 34 -4 37
rect 13 34 20 37
rect -30 20 -23 23
rect -19 20 1 23
rect -81 13 -75 16
rect -61 13 -53 16
rect -61 11 -58 13
rect -39 13 -22 16
rect -39 11 -36 13
rect -64 8 -58 11
rect -42 8 -36 11
rect -76 -3 -73 0
rect -54 -3 -51 0
rect -76 -6 -42 -3
<< m2contact >>
rect 60 5 68 11
rect -42 -7 -37 -2
<< pm12contact >>
rect 60 25 68 31
<< pdm12contact >>
rect 60 15 68 21
<< ndm12contact >>
rect -24 51 -19 56
rect 0 51 5 56
<< metal2 >>
rect -19 52 0 56
rect -24 47 -21 51
rect -8 50 -4 52
rect -33 44 -21 47
rect -33 -3 -30 44
rect -37 -6 -30 -3
<< labels >>
rlabel metal1 -74 65 -74 65 1 VDD
rlabel metal1 -54 72 -54 72 5 clk
rlabel metal1 -60 -5 -60 -5 1 gnd
rlabel pm12contact 64 28 64 28 7 poly_m1_m2
rlabel pdm12contact 63 18 63 18 7 pdiff_m1_m2
rlabel m2contact 63 8 63 8 7 m2contact
rlabel metal1 -79 14 -79 14 3 D
rlabel metal1 25 45 25 45 1 Q
<< end >>
