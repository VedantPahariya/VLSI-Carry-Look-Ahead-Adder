.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd

* Supply
Vdd vdd gnd 'SUPPLY'

* SPICE3 file created from complete.ext - technology: scmos

.option scale=0.09u

M1000 a_296_n76# clk a_278_n59# w_243_n62# CMOSP w=40 l=2
+  ad=160 pd=88 as=200 ps=90
M1001 gnd B_0 Pt0 Gnd CMOSN w=40 l=2
+  ad=6205 pd=3112 as=400 ps=180
M1002 VDD a_300_n163# a_296_n160# w_137_n171# CMOSP w=40 l=2
+  ad=11800 pd=5570 as=160 ps=88
M1003 a_44_n222# G0 gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1004 a_150_n274# C1 VDD w_137_n280# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1005 a_n101_n391# A_3 VDD w_n131_n463# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1006 a_198_n75# clk a_180_n58# w_123_n108# CMOSP w=40 l=2
+  ad=160 pd=88 as=200 ps=90
M1007 a_190_n274# a_174_n296# VDD w_137_n280# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1008 a_174_n405# a_150_n383# VDD w_137_n389# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1009 s_0 C0 pgxor0 w_38_n97# CMOSP w=8 l=2
+  ad=80 pd=52 as=120 ps=78
M1010 gnd a_278_n59# a_274_n24# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=80 ps=48
M1011 a_150_n165# C0 VDD w_137_n171# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1012 a_n30_n423# A_3 gnd Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1013 a_n101_n282# A_2 VDD w_n131_n354# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1014 a_190_n165# a_174_n187# VDD w_137_n171# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1015 a_149_n338# Cout VDD w_143_n351# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1016 C1 a_75_n113# VDD w_38_n97# CMOSP w=20 l=2
+  ad=160 pd=78 as=0 ps=0
M1017 a_174_n296# a_150_n274# VDD w_137_n280# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1018 a_44_n440# G2 a_51_n418# w_38_n424# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1019 a_n30_n314# A_2 gnd Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1020 a_195_n452# Pout gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1021 gnd a_254_n361# a_250_n326# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=80 ps=48
M1022 a_n101_n173# A_1 VDD w_n131_n245# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1023 gnd Pt3 P32 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1024 a_44_n222# G0 a_51_n200# w_38_n206# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1025 a_231_n296# C3 VDD w_137_n280# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1026 VDD G3 GPG3 w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1027 a_174_n187# a_150_n165# VDD w_137_n171# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1028 a_44_n331# G1 a_51_n309# w_38_n315# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1029 a_n30_n96# A_0 gnd Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1030 a_n30_n205# A_1 gnd Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1031 VDD G1 GPG1 w_38_n206# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1032 gnd a_254_n252# a_250_n217# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=80 ps=48
M1033 gnd Pt2 P21 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1034 gnd a_174_n296# a_183_n296# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1035 a_250_n326# clk Cout Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1036 a_231_n187# C2 VDD w_137_n171# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1037 VDD G2 GPG2 w_38_n315# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1038 gnd a_254_n143# a_250_n108# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=80 ps=48
M1039 a_150_n383# P32 a_150_n415# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1040 gnd Pt1 P10 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1041 gnd a_174_n187# a_183_n187# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1042 a_44_n440# G2 gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1043 a_174_n296# a_150_n274# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1044 a_n101_n64# A_0 VDD w_n131_n136# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1045 a_250_n217# clk S3 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1046 a_150_n165# P10 a_150_n197# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1047 a_174_n405# a_150_n383# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1048 VDD a_278_n59# a_254_n59# w_243_n62# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1049 a_274_n326# clk a_254_n361# Gnd CMOSN w=20 l=2
+  ad=80 pd=48 as=100 ps=50
M1050 a_231_n296# C3 gnd Gnd CMOSN w=10 l=2
+  ad=70 pd=48 as=0 ps=0
M1051 a_150_n274# P21 a_150_n306# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1052 VDD B_0 G0 w_n131_n136# CMOSP w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1053 a_250_n108# clk S2 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1054 a_174_n187# a_150_n165# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1055 pgxor1 C1 s_1 w_123_n108# CMOSP w=8 l=2
+  ad=125 pd=80 as=80 ps=52
M1056 VDD a_254_n361# Cout w_243_n364# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1057 a_231_n187# C2 gnd Gnd CMOSN w=10 l=2
+  ad=70 pd=48 as=0 ps=0
M1058 a_274_n217# clk a_254_n252# Gnd CMOSN w=20 l=2
+  ad=80 pd=48 as=100 ps=50
M1059 a_195_n452# Pout a_195_n460# w_189_n473# CMOSP w=40 l=2
+  ad=200 pd=90 as=240 ps=92
M1060 a_152_n23# clk S0 Gnd CMOSN w=20 l=2
+  ad=80 pd=48 as=100 ps=50
M1061 VDD S2 a_189_n117# w_205_n123# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1062 a_136_n124# C1 VDD w_123_n108# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1063 VDD a_254_n252# S3 w_137_n280# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1064 Gout GPG3 gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1065 a_51_n91# Pt0 VDD w_38_n97# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1066 a_274_n108# clk a_254_n143# Gnd CMOSN w=20 l=2
+  ad=80 pd=48 as=100 ps=50
M1067 pgxor0 B_0 a_n101_n64# Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=70 ps=48
M1068 VDD G0 C1 w_38_n97# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1069 pgxor1 a_136_n124# s_1 Gnd CMOSN w=4 l=2
+  ad=69 pd=58 as=40 ps=36
M1070 VDD a_254_n143# S2 w_137_n171# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1071 gnd C4 a_300_n381# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1072 VDD P32 a_150_n383# w_137_n389# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1073 a_91_n341# a_75_n331# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1074 C4 a_216_n386# a_257_n392# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1075 gnd a_180_n58# a_176_n23# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=80 ps=48
M1076 a_136_n124# C1 gnd Gnd CMOSN w=10 l=2
+  ad=70 pd=48 as=0 ps=0
M1077 VDD s_1 a_318_n76# w_243_n62# CMOSP w=40 l=2
+  ad=0 pd=0 as=160 ps=88
M1078 a_91_n232# a_75_n222# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1079 gnd s_3 a_300_n272# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1080 pgxor0 B_0 A_0 w_n47_n53# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1081 VDD P21 a_150_n274# w_137_n280# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 gnd Pt0 a_44_n123# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1083 P32 Pt2 a_76_n374# w_38_n424# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1084 a_183_n296# GPG2 a_190_n274# w_137_n280# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1085 gnd C0bar a_195_n452# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1086 VDD a_216_n386# C4 w_137_n389# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1087 VDD s_0 a_220_n75# w_123_n108# CMOSP w=40 l=2
+  ad=0 pd=0 as=160 ps=88
M1088 a_91_n123# a_75_n113# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1089 gnd s_2 a_300_n163# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1090 VDD P10 a_150_n165# w_137_n171# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 gnd a_300_n381# a_278_n361# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1092 gnd a_278_n361# a_274_n326# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1093 P21 Pt1 a_76_n265# w_38_n315# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1094 a_183_n187# GPG1 a_190_n165# w_137_n171# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1095 gnd a_278_n252# a_274_n217# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 C3 a_183_n296# VDD w_137_n280# CMOSP w=20 l=2
+  ad=140 pd=76 as=0 ps=0
M1097 gnd a_300_n272# a_278_n252# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1098 pgxor2 B_2 a_n101_n282# Gnd CMOSN w=4 l=2
+  ad=69 pd=58 as=70 ps=48
M1099 P10 Pt0 a_76_n156# w_38_n206# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1100 VDD a_300_n79# a_296_n76# w_243_n62# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 gnd a_278_n143# a_274_n108# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 C2 a_183_n187# VDD w_137_n171# CMOSP w=20 l=2
+  ad=140 pd=76 as=0 ps=0
M1103 pgxor3 B_3 A_3 w_n47_n380# CMOSP w=8 l=2
+  ad=125 pd=80 as=40 ps=26
M1104 VDD a_180_n58# a_156_n58# w_123_n108# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1105 gnd a_300_n163# a_278_n143# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1106 pgxor1 B_1 a_n101_n173# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=70 ps=48
M1107 Gout GPG3 a_198_n403# w_137_n389# CMOSP w=40 l=2
+  ad=200 pd=90 as=240 ps=92
M1108 a_183_n296# GPG2 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 a_44_n123# C0bar a_51_n91# w_38_n97# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1110 C0 a_84_n59# s_0 Gnd CMOSN w=4 l=2
+  ad=29 pd=22 as=40 ps=36
M1111 pgxor2 a_231_n187# s_2 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1112 VDD a_202_n78# a_198_n75# w_123_n108# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 G0 A_0 VDD w_n131_n136# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 a_183_n187# GPG1 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 pgxor2 B_2 A_2 w_n47_n271# CMOSP w=8 l=2
+  ad=125 pd=80 as=40 ps=26
M1116 VDD S1 a_333_n98# w_243_n62# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1117 pgxor3 C3 s_3 w_137_n280# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=52
M1118 a_216_n386# a_195_n452# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1119 a_216_n386# a_195_n452# VDD w_189_n473# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1120 a_91_n450# a_75_n440# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1121 C3 a_183_n296# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1122 a_195_n460# C0bar VDD w_189_n473# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 VDD A_3 a_n125_n450# w_n131_n463# CMOSP w=80 l=2
+  ad=0 pd=0 as=480 ps=172
M1124 VDD a_278_n361# a_254_n361# w_243_n364# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1125 C0 pgxor0 s_0 w_38_n97# CMOSP w=8 l=2
+  ad=45 pd=28 as=0 ps=0
M1126 gnd S2 a_189_n117# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1127 pgxor1 B_1 A_1 w_n47_n162# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1128 pgxor2 C2 s_2 w_137_n171# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=52
M1129 VDD B_3 G3 w_n131_n463# CMOSP w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1130 C0bar C0 VDD w_n131_n136# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1131 C2 a_183_n187# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1132 gnd a_174_n405# Gout Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 VDD A_2 a_n125_n341# w_n131_n354# CMOSP w=80 l=2
+  ad=0 pd=0 as=480 ps=172
M1134 a_274_n24# clk a_254_n59# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1135 VDD a_278_n252# a_254_n252# w_137_n280# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1136 s_1 pgxor1 a_136_n124# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1137 VDD B_1 G1 w_n131_n245# CMOSP w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1138 Pt3 A_3 gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1139 VDD B_2 G2 w_n131_n354# CMOSP w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1140 gnd S1 a_333_n98# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1141 VDD S0 a_153_n133# w_137_n171# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1142 gnd S0 a_153_n133# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1143 VDD A_1 a_n125_n232# w_n131_n245# CMOSP w=80 l=2
+  ad=0 pd=0 as=480 ps=172
M1144 a_149_n229# S3 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1145 gnd Pt2 a_44_n331# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1146 a_176_n23# clk a_156_n58# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1147 VDD a_278_n143# a_254_n143# w_137_n171# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1148 gnd P10 a_156_n444# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1149 Pt2 A_2 gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1150 a_318_n76# clk a_300_n79# w_243_n62# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1151 a_296_n378# clk a_278_n361# w_243_n364# CMOSP w=40 l=2
+  ad=160 pd=88 as=200 ps=90
M1152 gnd Pt1 a_44_n222# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 a_257_n392# Gout gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 VDD A_0 a_n125_n123# w_n131_n136# CMOSP w=80 l=2
+  ad=0 pd=0 as=480 ps=172
M1155 pgxor3 B_3 a_n101_n391# Gnd CMOSN w=4 l=2
+  ad=69 pd=58 as=70 ps=48
M1156 C0bar C0 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1157 Pt1 A_1 gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1158 gnd a_254_n59# a_250_n24# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=80 ps=48
M1159 a_220_n75# clk a_202_n78# w_123_n108# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1160 a_296_n269# clk a_278_n252# w_137_n280# CMOSP w=40 l=2
+  ad=160 pd=88 as=200 ps=90
M1161 VDD P10 Pout w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1162 a_75_n331# a_44_n331# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1163 GPG2 G2 a_91_n341# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1164 a_76_n374# Pt3 VDD w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 Pt0 A_0 gnd Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 C4 Gout VDD w_137_n389# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 pgxor3 a_231_n296# s_3 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1168 gnd a_156_n58# a_152_n23# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1169 a_n101_n64# A_0 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 a_296_n160# clk a_278_n143# w_137_n171# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1171 a_75_n222# a_44_n222# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1172 GPG1 G1 a_91_n232# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1173 a_51_n418# Pt3 VDD w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1174 a_44_n123# C0bar gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 a_76_n265# Pt2 VDD w_38_n315# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 B_2 a_n101_n282# pgxor2 Gnd CMOSN w=4 l=2
+  ad=29 pd=22 as=0 ps=0
M1177 a_51_n200# Pt1 VDD w_38_n206# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 G3 B_3 a_n30_n423# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1179 a_75_n113# a_44_n123# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1180 GPG3 a_75_n440# VDD w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 C1 G0 a_91_n123# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1182 a_76_n156# Pt1 VDD w_38_n206# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 a_51_n309# Pt2 VDD w_38_n315# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1184 G1 B_1 a_n30_n205# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1185 B_3 A_3 pgxor3 w_n47_n380# CMOSP w=8 l=2
+  ad=45 pd=28 as=0 ps=0
M1186 B_1 a_n101_n173# pgxor1 Gnd CMOSN w=4 l=2
+  ad=29 pd=22 as=0 ps=0
M1187 GPG1 a_75_n222# VDD w_38_n206# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 G2 B_2 a_n30_n314# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1189 s_2 pgxor2 a_231_n187# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 a_75_n440# a_44_n440# VDD w_38_n424# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1191 GPG2 a_75_n331# VDD w_38_n315# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 a_198_n403# a_174_n405# VDD w_137_n389# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1193 P32 Pt2 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 s_1 pgxor1 C1 w_123_n108# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 VDD a_254_n59# S1 w_243_n62# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1196 B_2 A_2 pgxor2 w_n47_n271# CMOSP w=8 l=2
+  ad=45 pd=28 as=0 ps=0
M1197 a_150_n415# GPG1 gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 G0 B_0 a_n30_n96# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1199 a_75_n222# a_44_n222# VDD w_38_n206# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1200 s_3 pgxor3 C3 w_137_n280# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1201 gnd Pt3 a_44_n440# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1202 a_149_n338# Cout gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1203 P21 Pt1 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1204 a_75_n331# a_44_n331# VDD w_38_n315# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1205 a_150_n197# C0 gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1206 gnd s_1 a_300_n79# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1207 a_150_n306# C1 gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 VDD a_156_n58# S0 w_123_n108# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1209 B_1 A_1 pgxor1 w_n47_n162# CMOSP w=8 l=2
+  ad=45 pd=28 as=0 ps=0
M1210 a_n125_n450# B_3 Pt3 w_n131_n463# CMOSP w=80 l=2
+  ad=0 pd=0 as=400 ps=170
M1211 VDD C4 a_318_n378# w_243_n364# CMOSP w=40 l=2
+  ad=0 pd=0 as=160 ps=88
M1212 s_2 pgxor2 C2 w_137_n171# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1213 P10 Pt0 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 a_n101_n391# A_3 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 a_149_n229# S3 VDD w_143_n242# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1216 G3 A_3 VDD w_n131_n463# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 gnd s_0 a_202_n78# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1218 B_0 a_n101_n64# pgxor0 Gnd CMOSN w=4 l=2
+  ad=29 pd=22 as=0 ps=0
M1219 a_75_n440# a_44_n440# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1220 a_84_n59# pgxor0 VDD w_38_n97# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1221 VDD s_3 a_318_n269# w_137_n280# CMOSP w=40 l=2
+  ad=0 pd=0 as=160 ps=88
M1222 GPG3 G3 a_91_n450# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1223 a_n125_n341# B_2 Pt2 w_n131_n354# CMOSP w=80 l=2
+  ad=0 pd=0 as=400 ps=170
M1224 gnd B_3 Pt3 Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 a_318_n378# clk a_300_n381# w_243_n364# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1226 G2 A_2 VDD w_n131_n354# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 a_n101_n282# A_2 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 a_75_n113# a_44_n123# VDD w_38_n97# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1229 a_n125_n232# B_1 Pt1 w_n131_n245# CMOSP w=80 l=2
+  ad=0 pd=0 as=400 ps=170
M1230 VDD s_2 a_318_n160# w_137_n171# CMOSP w=40 l=2
+  ad=0 pd=0 as=160 ps=88
M1231 a_156_n444# P32 Pout Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1232 a_318_n269# clk a_300_n272# w_137_n280# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1233 VDD a_300_n381# a_296_n378# w_243_n364# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1234 gnd B_2 Pt2 Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 a_n101_n173# A_1 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1236 G1 A_1 VDD w_n131_n245# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1237 B_3 a_n101_n391# pgxor3 Gnd CMOSN w=4 l=2
+  ad=29 pd=22 as=0 ps=0
M1238 a_250_n24# clk S1 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1239 gnd a_300_n79# a_278_n59# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1240 B_0 A_0 pgxor0 w_n47_n53# CMOSP w=8 l=2
+  ad=45 pd=28 as=0 ps=0
M1241 a_n125_n123# B_0 Pt0 w_n131_n136# CMOSP w=80 l=2
+  ad=0 pd=0 as=400 ps=170
M1242 a_44_n331# G1 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1243 a_84_n59# pgxor0 gnd Gnd CMOSN w=10 l=2
+  ad=70 pd=48 as=0 ps=0
M1244 a_318_n160# clk a_300_n163# w_137_n171# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1245 gnd B_1 Pt1 Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1246 VDD a_300_n272# a_296_n269# w_137_n280# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1247 a_150_n383# GPG1 VDD w_137_n389# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1248 s_0 C0 a_84_n59# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1249 Pout P32 VDD w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1250 gnd a_202_n78# a_180_n58# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1251 s_3 pgxor3 a_231_n296# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_300_n381# C4 0.05fF
C1 G2 a_44_n440# 0.06fF
C2 a_202_n78# s_0 0.05fF
C3 pgxor2 VDD 0.24fF
C4 A_0 VDD 0.81fF
C5 S3 w_137_n280# 0.14fF
C6 a_174_n405# GPG3 0.14fF
C7 P32 Pt3 0.14fF
C8 A_3 a_n101_n391# 0.12fF
C9 s_2 a_231_n187# 0.12fF
C10 B_3 C0bar 0.00fF
C11 clk S2 0.19fF
C12 S3 a_300_n272# 0.12fF
C13 a_75_n222# gnd 0.06fF
C14 B_1 a_n101_n173# 0.20fF
C15 a_n101_n64# w_n131_n136# 0.02fF
C16 G0 w_38_n97# 0.06fF
C17 Pt3 C0bar 0.00fF
C18 S2 VDD 0.78fF
C19 G1 VDD 0.33fF
C20 P21 a_150_n274# 0.06fF
C21 s_3 C3 0.10fF
C22 pgxor1 gnd 0.99fF
C23 s_1 gnd 0.44fF
C24 a_n101_n64# pgxor0 0.12fF
C25 C3 pgxor3 0.22fF
C26 s_3 gnd 0.02fF
C27 w_38_n97# C1 0.05fF
C28 pgxor1 C0 0.06fF
C29 Pt0 VDD 0.21fF
C30 GPG2 gnd 0.04fF
C31 a_75_n440# G3 0.09fF
C32 B_2 G2 0.37fF
C33 pgxor3 gnd 0.90fF
C34 a_183_n296# VDD 0.03fF
C35 a_n101_n64# B_0 0.20fF
C36 G0 C0bar 0.02fF
C37 Pt2 a_44_n331# 0.09fF
C38 GPG1 C1 0.29fF
C39 Gout a_216_n386# 0.31fF
C40 s_0 pgxor0 0.10fF
C41 a_296_n269# VDD 0.01fF
C42 VDD w_137_n389# 0.28fF
C43 clk VDD 0.95fF
C44 a_44_n331# w_38_n315# 0.10fF
C45 GPG1 a_183_n187# 0.23fF
C46 a_202_n78# w_123_n108# 0.09fF
C47 G2 gnd 1.26fF
C48 G0 A_0 0.16fF
C49 B_1 w_n131_n245# 0.44fF
C50 P10 gnd 0.56fF
C51 pgxor1 a_136_n124# 0.05fF
C52 s_1 a_136_n124# 0.12fF
C53 s_0 S0 0.07fF
C54 C4 w_243_n364# 0.20fF
C55 w_n131_n463# gnd 0.03fF
C56 pgxor3 A_3 0.11fF
C57 a_300_n79# S1 0.12fF
C58 P10 C0 0.32fF
C59 a_150_n165# VDD 0.02fF
C60 a_250_n108# gnd 0.01fF
C61 pgxor3 a_n101_n391# 0.12fF
C62 a_149_n338# gnd 0.07fF
C63 a_195_n452# Pout 0.22fF
C64 s_0 a_84_n59# 0.12fF
C65 pgxor2 C1 0.36fF
C66 B_3 VDD 0.06fF
C67 Pt3 VDD 0.14fF
C68 G0 Pt0 0.88fF
C69 a_n125_n341# C0bar 0.00fF
C70 GPG1 GPG3 0.00fF
C71 Pt1 gnd 0.43fF
C72 A_3 w_n131_n463# 0.48fF
C73 A_1 C0bar 0.00fF
C74 Cout a_149_n338# 0.04fF
C75 a_216_n386# gnd 0.05fF
C76 a_51_n418# VDD 0.01fF
C77 a_n101_n391# w_n131_n463# 0.02fF
C78 S0 a_220_n75# 0.00fF
C79 a_300_n163# gnd 0.04fF
C80 a_195_n452# w_189_n473# 0.10fF
C81 B_3 Pt3 0.20fF
C82 a_150_n383# a_174_n405# 0.04fF
C83 P32 GPG3 0.17fF
C84 a_n101_n64# gnd 0.28fF
C85 pgxor1 s_1 0.52fF
C86 a_189_n117# w_205_n123# 0.02fF
C87 a_153_n133# w_137_n171# 0.02fF
C88 a_156_n444# gnd 0.02fF
C89 G0 VDD 0.29fF
C90 a_183_n296# w_137_n280# 0.10fF
C91 a_300_n163# s_2 0.05fF
C92 a_278_n252# clk 0.33fF
C93 a_254_n252# gnd 0.08fF
C94 B_3 w_n47_n380# 0.28fF
C95 a_44_n222# VDD 0.08fF
C96 w_137_n171# a_254_n143# 0.11fF
C97 S0 w_123_n108# 0.43fF
C98 a_195_n460# VDD 0.02fF
C99 a_278_n252# VDD 0.08fF
C100 A_2 Pt2 0.09fF
C101 s_3 pgxor3 0.54fF
C102 a_174_n296# a_183_n296# 0.13fF
C103 w_143_n242# gnd 0.04fF
C104 w_243_n62# clk 0.37fF
C105 s_0 gnd 0.30fF
C106 w_137_n280# clk 0.37fF
C107 a_174_n405# Gout 0.09fF
C108 a_333_n98# gnd 0.02fF
C109 A_1 G1 0.16fF
C110 a_274_n217# gnd 0.01fF
C111 a_300_n272# clk 0.03fF
C112 w_243_n62# VDD 0.14fF
C113 w_137_n280# VDD 0.36fF
C114 a_300_n79# gnd 0.04fF
C115 s_0 C0 0.57fF
C116 C0bar w_n47_n53# 0.38fF
C117 C1 VDD 0.22fF
C118 a_150_n274# gnd 0.04fF
C119 S1 a_278_n59# 0.12fF
C120 a_44_n440# a_75_n440# 0.04fF
C121 a_300_n272# VDD 0.08fF
C122 S0 w_137_n171# 0.11fF
C123 a_231_n296# clk 0.19fF
C124 P32 Pout 0.15fF
C125 a_174_n296# VDD 0.02fF
C126 a_183_n187# VDD 0.03fF
C127 GPG2 G2 0.06fF
C128 P10 pgxor1 0.29fF
C129 Pout C0bar 0.08fF
C130 pgxor3 G2 0.75fF
C131 A_0 w_n47_n53# 0.19fF
C132 A_2 w_n131_n354# 0.48fF
C133 a_254_n361# w_243_n364# 0.11fF
C134 P10 GPG2 0.05fF
C135 GPG1 P21 0.04fF
C136 G2 w_38_n424# 0.22fF
C137 GPG1 w_38_n206# 0.21fF
C138 a_44_n331# gnd 0.12fF
C139 P10 pgxor3 0.05fF
C140 a_278_n361# gnd 0.06fF
C141 a_n101_n282# w_n131_n354# 0.02fF
C142 P10 w_38_n424# 0.17fF
C143 a_75_n331# VDD 0.08fF
C144 B_1 gnd 0.11fF
C145 S2 w_205_n123# 0.10fF
C146 Pt2 P32 0.28fF
C147 A_1 VDD 0.28fF
C148 gnd a_278_n143# 0.06fF
C149 C4 w_137_n389# 0.05fF
C150 a_44_n222# G0 0.06fF
C151 a_300_n381# gnd 0.04fF
C152 C4 clk 0.61fF
C153 Pt2 C0bar 0.00fF
C154 w_38_n97# pgxor0 0.31fF
C155 GPG3 w_137_n389# 0.50fF
C156 w_189_n473# C0bar 0.18fF
C157 a_174_n405# gnd 0.06fF
C158 a_156_n58# w_123_n108# 0.11fF
C159 C4 VDD 0.08fF
C160 w_n131_n245# C0bar 0.20fF
C161 a_278_n361# Cout 0.12fF
C162 GPG3 VDD 0.07fF
C163 pgxor2 P21 0.45fF
C164 a_250_n24# gnd 0.01fF
C165 w_n47_n162# pgxor1 0.07fF
C166 G0 C1 0.06fF
C167 a_152_n23# gnd 0.01fF
C168 w_n131_n136# C0bar 0.30fF
C169 G0 a_n30_n96# 0.02fF
C170 GPG1 a_150_n383# 0.04fF
C171 a_278_n252# w_137_n280# 0.12fF
C172 C2 gnd 0.02fF
C173 Cout a_300_n381# 0.12fF
C174 a_n125_n123# C0bar 0.00fF
C175 w_137_n171# gnd 0.06fF
C176 a_278_n59# gnd 0.06fF
C177 G3 VDD 0.12fF
C178 w_n131_n354# C0bar 0.20fF
C179 G1 w_38_n206# 0.06fF
C180 a_318_n378# VDD 0.01fF
C181 G1 Pt2 0.20fF
C182 w_137_n171# C0 0.12fF
C183 w_205_n123# VDD 0.03fF
C184 pgxor0 C0bar 0.51fF
C185 P32 a_150_n383# 0.06fF
C186 w_137_n280# C1 0.12fF
C187 w_38_n97# a_84_n59# 0.02fF
C188 w_n131_n136# A_0 0.49fF
C189 s_2 C2 0.10fF
C190 a_333_n98# s_1 0.02fF
C191 a_300_n272# w_137_n280# 0.09fF
C192 a_180_n58# S0 0.12fF
C193 s_2 w_137_n171# 0.28fF
C194 a_195_n452# gnd 0.18fF
C195 G1 w_n131_n245# 0.06fF
C196 P10 Pt1 0.14fF
C197 a_300_n79# s_1 0.05fF
C198 G1 w_38_n315# 0.22fF
C199 a_174_n296# w_137_n280# 0.14fF
C200 a_136_n124# w_123_n108# 0.03fF
C201 a_174_n187# w_137_n171# 0.14fF
C202 w_38_n206# Pt0 0.14fF
C203 Pout VDD 0.14fF
C204 a_231_n296# w_137_n280# 0.02fF
C205 B_2 A_2 0.32fF
C206 C0bar B_0 0.02fF
C207 pgxor0 A_0 0.11fF
C208 B_3 G3 0.37fF
C209 Cout a_296_n378# 0.01fF
C210 a_44_n123# a_75_n113# 0.04fF
C211 S1 a_296_n76# 0.01fF
C212 a_150_n274# GPG2 0.07fF
C213 S3 a_318_n269# 0.01fF
C214 a_202_n78# clk 0.03fF
C215 Pt3 G3 0.77fF
C216 B_2 a_n101_n282# 0.20fF
C217 S3 gnd 0.15fF
C218 a_202_n78# VDD 0.08fF
C219 S2 a_254_n143# 0.17fF
C220 a_318_n76# VDD 0.01fF
C221 A_2 gnd 0.07fF
C222 gnd a_75_n113# 0.06fF
C223 A_0 B_0 0.32fF
C224 w_n131_n136# Pt0 0.04fF
C225 P21 VDD 0.32fF
C226 C0 a_75_n113# 0.00fF
C227 w_38_n97# a_44_n123# 0.09fF
C228 B_1 pgxor1 0.52fF
C229 w_38_n206# VDD 0.16fF
C230 a_n101_n282# gnd 0.28fF
C231 Pt2 VDD 0.25fF
C232 C2 a_231_n187# 0.23fF
C233 w_189_n473# VDD 0.07fF
C234 a_231_n187# w_137_n171# 0.02fF
C235 B_2 w_n47_n271# 0.28fF
C236 gnd a_176_n23# 0.01fF
C237 Cout w_143_n351# 0.06fF
C238 w_n131_n245# VDD 0.18fF
C239 S2 S0 0.00fF
C240 w_38_n315# VDD 0.16fF
C241 w_38_n97# gnd 0.10fF
C242 a_150_n306# gnd 0.02fF
C243 a_254_n361# clk 0.09fF
C244 pgxor1 w_123_n108# 0.41fF
C245 s_1 w_123_n108# 0.14fF
C246 a_189_n117# gnd 0.13fF
C247 w_38_n97# C0 0.95fF
C248 w_n131_n136# VDD 0.24fF
C249 a_296_n160# S2 0.01fF
C250 a_254_n361# VDD 0.09fF
C251 Cout w_243_n364# 0.14fF
C252 Pt0 B_0 0.20fF
C253 GPG1 gnd 0.18fF
C254 a_153_n133# VDD 0.15fF
C255 clk a_254_n143# 0.09fF
C256 a_198_n75# VDD 0.01fF
C257 B_2 C0bar 0.00fF
C258 a_180_n58# gnd 0.06fF
C259 C0bar a_44_n123# 0.06fF
C260 w_n131_n354# VDD 0.18fF
C261 Pt2 Pt3 0.07fF
C262 GPG1 C0 0.04fF
C263 a_250_n326# gnd 0.01fF
C264 VDD a_254_n143# 0.09fF
C265 pgxor0 VDD 1.00fF
C266 a_150_n383# w_137_n389# 0.15fF
C267 P32 gnd 0.32fF
C268 Pout a_195_n460# 0.04fF
C269 G1 a_n30_n205# 0.02fF
C270 a_174_n187# GPG1 0.14fF
C271 a_150_n383# VDD 0.02fF
C272 C0bar gnd 0.47fF
C273 pgxor2 B_2 0.52fF
C274 clk S1 0.19fF
C275 clk S0 0.21fF
C276 a_75_n440# w_38_n424# 0.10fF
C277 B_0 VDD 0.06fF
C278 C0bar C0 0.06fF
C279 S1 VDD 0.64fF
C280 S0 VDD 0.70fF
C281 Gout w_137_n389# 0.23fF
C282 G0 w_38_n206# 0.22fF
C283 clk a_254_n59# 0.09fF
C284 a_44_n440# VDD 0.08fF
C285 A_0 gnd 0.07fF
C286 pgxor2 gnd 1.03fF
C287 a_44_n222# w_38_n206# 0.10fF
C288 Gout VDD 0.12fF
C289 a_254_n59# VDD 0.09fF
C290 a_84_n59# VDD 0.21fF
C291 a_296_n160# VDD 0.01fF
C292 B_1 Pt1 0.20fF
C293 s_2 pgxor2 0.54fF
C294 A_3 C0bar 0.00fF
C295 S2 gnd 0.09fF
C296 P21 w_137_n280# 0.06fF
C297 S3 s_3 0.06fF
C298 P10 w_137_n171# 0.06fF
C299 G1 gnd 1.26fF
C300 P21 C1 0.09fF
C301 Pt0 a_44_n123# 0.09fF
C302 A_1 a_n101_n173# 0.12fF
C303 G0 w_n131_n136# 0.06fF
C304 B_1 w_n47_n162# 0.28fF
C305 GPG3 G3 0.06fF
C306 s_2 S2 0.06fF
C307 Pt3 a_44_n440# 0.09fF
C308 a_183_n296# C3 0.04fF
C309 Pt0 gnd 0.28fF
C310 a_149_n229# gnd 0.07fF
C311 a_n125_n450# C0bar 0.00fF
C312 Pt0 C0 0.01fF
C313 a_183_n296# gnd 0.12fF
C314 B_2 VDD 0.06fF
C315 VDD a_44_n123# 0.04fF
C316 A_2 G2 0.16fF
C317 C3 VDD 0.09fF
C318 G0 B_0 0.37fF
C319 clk gnd 2.84fF
C320 clk a_156_n58# 0.09fF
C321 a_318_n269# VDD 0.01fF
C322 a_231_n187# pgxor2 0.16fF
C323 a_n125_n232# C0bar 0.00fF
C324 a_149_n338# w_143_n351# 0.02fF
C325 GPG1 GPG2 0.05fF
C326 VDD gnd 1.64fF
C327 a_300_n163# w_137_n171# 0.09fF
C328 a_75_n331# w_38_n315# 0.10fF
C329 a_156_n58# VDD 0.09fF
C330 s_0 w_123_n108# 0.24fF
C331 GPG1 pgxor3 0.05fF
C332 s_2 clk 0.61fF
C333 A_1 w_n131_n245# 0.48fF
C334 VDD C0 3.15fF
C335 a_216_n386# a_195_n452# 0.04fF
C336 w_243_n62# S1 0.21fF
C337 a_51_n309# VDD 0.01fF
C338 a_150_n165# gnd 0.04fF
C339 s_2 VDD 0.06fF
C340 pgxor3 P32 0.46fF
C341 Cout clk 0.19fF
C342 a_91_n341# gnd 0.02fF
C343 a_174_n187# VDD 0.02fF
C344 a_150_n165# C0 0.04fF
C345 P32 w_38_n424# 0.19fF
C346 B_3 gnd 0.11fF
C347 w_243_n62# a_254_n59# 0.11fF
C348 Cout VDD 1.23fF
C349 a_75_n222# G1 0.09fF
C350 Pt3 gnd 0.60fF
C351 P10 GPG1 0.50fF
C352 a_150_n165# a_174_n187# 0.04fF
C353 A_3 VDD 0.28fF
C354 P10 P32 0.46fF
C355 a_254_n252# S3 0.17fF
C356 a_231_n187# clk 0.19fF
C357 a_n101_n173# w_n131_n245# 0.02fF
C358 B_3 A_3 0.32fF
C359 C0bar w_n131_n463# 0.20fF
C360 Pout w_189_n473# 0.26fF
C361 S3 w_143_n242# 0.06fF
C362 B_3 a_n101_n391# 0.20fF
C363 a_150_n383# GPG3 0.07fF
C364 A_3 Pt3 0.09fF
C365 G0 gnd 1.58fF
C366 pgxor1 Pt0 0.27fF
C367 a_44_n222# gnd 0.12fF
C368 P10 pgxor2 0.08fF
C369 G0 C0 0.35fF
C370 C3 w_137_n280# 0.27fF
C371 a_278_n252# gnd 0.06fF
C372 A_3 w_n47_n380# 0.19fF
C373 a_75_n222# VDD 0.08fF
C374 w_137_n171# a_278_n143# 0.12fF
C375 pgxor0 w_n47_n53# 0.07fF
C376 C4 Gout 0.02fF
C377 a_274_n108# gnd 0.01fF
C378 GPG2 a_183_n296# 0.23fF
C379 P21 Pt2 0.14fF
C380 GPG3 Gout 0.22fF
C381 clk pgxor1 0.06fF
C382 C1 gnd 0.34fF
C383 clk s_1 1.61fF
C384 C3 a_231_n296# 0.23fF
C385 a_300_n272# gnd 0.04fF
C386 s_3 clk 0.61fF
C387 Pt1 C0bar 0.00fF
C388 w_38_n97# s_0 0.07fF
C389 P21 w_38_n315# 0.08fF
C390 pgxor1 VDD 0.25fF
C391 C1 C0 0.11fF
C392 B_0 w_n47_n53# 0.28fF
C393 s_1 VDD 0.06fF
C394 a_174_n296# gnd 0.02fF
C395 a_183_n187# gnd 0.12fF
C396 s_3 VDD 0.06fF
C397 VDD a_51_n91# 0.01fF
C398 Pt2 w_38_n315# 0.25fF
C399 GPG2 VDD 0.04fF
C400 P10 Pt0 0.28fF
C401 C2 w_137_n171# 0.27fF
C402 pgxor3 VDD 0.24fF
C403 Pt1 pgxor2 0.27fF
C404 VDD w_38_n424# 0.26fF
C405 a_278_n361# w_243_n364# 0.12fF
C406 a_174_n187# a_183_n187# 0.13fF
C407 a_75_n331# gnd 0.06fF
C408 Pt2 w_n131_n354# 0.04fF
C409 a_n101_n64# A_0 0.12fF
C410 P10 w_137_n389# 0.02fF
C411 G2 VDD 0.33fF
C412 Pt1 G1 0.85fF
C413 A_1 gnd 0.07fF
C414 a_318_n76# S1 0.01fF
C415 C1 a_136_n124# 0.09fF
C416 G2 a_n30_n314# 0.02fF
C417 a_202_n78# S0 0.08fF
C418 a_300_n381# w_243_n364# 0.09fF
C419 a_300_n163# S2 0.12fF
C420 pgxor3 B_3 0.52fF
C421 P10 VDD 0.19fF
C422 w_n131_n463# VDD 0.18fF
C423 C4 gnd 0.02fF
C424 Pt3 w_38_n424# 0.25fF
C425 a_44_n222# a_75_n222# 0.04fF
C426 Pt1 Pt0 0.07fF
C427 P10 a_150_n165# 0.06fF
C428 pgxor3 w_n47_n380# 0.07fF
C429 G2 Pt3 0.20fF
C430 G0 pgxor1 0.75fF
C431 w_n131_n136# B_0 0.44fF
C432 G3 gnd 1.04fF
C433 B_3 w_n131_n463# 0.44fF
C434 a_216_n386# w_137_n389# 0.08fF
C435 Cout C4 0.06fF
C436 B_1 C0bar 0.00fF
C437 w_205_n123# gnd 0.05fF
C438 a_180_n58# w_123_n108# 0.12fF
C439 Pt3 w_n131_n463# 0.04fF
C440 a_n101_n173# gnd 0.28fF
C441 a_153_n133# S0 0.05fF
C442 S0 a_198_n75# 0.01fF
C443 Pt1 VDD 0.25fF
C444 a_300_n163# clk 0.03fF
C445 a_216_n386# VDD 0.06fF
C446 pgxor0 B_0 0.52fF
C447 w_243_n62# s_1 0.20fF
C448 C1 pgxor1 0.77fF
C449 C1 s_1 0.11fF
C450 a_300_n163# VDD 0.08fF
C451 a_149_n229# w_143_n242# 0.02fF
C452 s_3 w_137_n280# 0.28fF
C453 Pout gnd 0.19fF
C454 a_n101_n64# VDD 0.02fF
C455 GPG2 w_137_n280# 0.35fF
C456 a_300_n272# s_3 0.05fF
C457 GPG1 w_137_n171# 0.35fF
C458 a_150_n197# gnd 0.02fF
C459 a_254_n252# clk 0.09fF
C460 GPG2 C1 0.02fF
C461 G1 a_44_n331# 0.06fF
C462 pgxor3 w_137_n280# 0.37fF
C463 Cout a_318_n378# 0.01fF
C464 pgxor0 a_84_n59# 0.23fF
C465 A_3 G3 0.16fF
C466 a_254_n252# VDD 0.09fF
C467 a_174_n296# GPG2 0.14fF
C468 s_3 a_231_n296# 0.12fF
C469 B_2 Pt2 0.20fF
C470 a_202_n78# gnd 0.04fF
C471 s_0 clk 0.73fF
C472 B_1 G1 0.37fF
C473 A_2 a_n101_n282# 0.12fF
C474 a_250_n217# gnd 0.01fF
C475 w_143_n242# VDD 0.02fF
C476 a_274_n24# gnd 0.01fF
C477 s_0 VDD 0.41fF
C478 clk a_300_n79# 0.03fF
C479 S2 a_278_n143# 0.12fF
C480 a_333_n98# VDD 0.02fF
C481 a_231_n296# pgxor3 0.16fF
C482 P21 gnd 0.29fF
C483 S1 a_254_n59# 0.17fF
C484 a_300_n79# VDD 0.08fF
C485 Pt2 gnd 0.43fF
C486 a_150_n274# VDD 0.02fF
C487 P10 w_137_n280# 0.02fF
C488 w_38_n97# a_75_n113# 0.10fF
C489 w_189_n473# gnd 0.10fF
C490 P10 C1 0.08fF
C491 A_1 pgxor1 0.11fF
C492 w_n131_n245# gnd 0.03fF
C493 C2 pgxor2 0.22fF
C494 a_195_n452# C0bar 0.10fF
C495 pgxor2 w_137_n171# 0.37fF
C496 B_2 w_n131_n354# 0.44fF
C497 A_2 w_n47_n271# 0.19fF
C498 a_91_n123# gnd 0.02fF
C499 w_n131_n136# gnd 0.14fF
C500 Pt1 G0 0.20fF
C501 a_91_n123# C0 0.00fF
C502 a_278_n361# clk 0.33fF
C503 a_254_n361# gnd 0.08fF
C504 a_44_n331# VDD 0.08fF
C505 Pt1 a_44_n222# 0.09fF
C506 a_n125_n123# gnd 0.01fF
C507 w_n131_n136# C0 0.13fF
C508 a_75_n331# G2 0.09fF
C509 S2 w_137_n171# 0.14fF
C510 a_318_n160# S2 0.01fF
C511 w_n131_n354# gnd 0.03fF
C512 a_278_n361# VDD 0.08fF
C513 B_1 VDD 0.06fF
C514 gnd a_254_n143# 0.08fF
C515 clk a_278_n143# 0.33fF
C516 A_2 C0bar 0.00fF
C517 a_220_n75# VDD 0.01fF
C518 pgxor0 gnd 0.02fF
C519 a_274_n326# gnd 0.01fF
C520 a_300_n381# clk 0.03fF
C521 VDD a_278_n143# 0.08fF
C522 pgxor0 C0 0.29fF
C523 GPG3 w_38_n424# 0.30fF
C524 a_174_n405# w_137_n389# 0.22fF
C525 clk w_123_n108# 0.44fF
C526 a_150_n383# gnd 0.04fF
C527 a_300_n381# VDD 0.08fF
C528 a_n101_n173# pgxor1 0.12fF
C529 a_254_n361# Cout 0.17fF
C530 a_174_n405# VDD 0.02fF
C531 B_0 gnd 0.12fF
C532 w_123_n108# VDD 0.16fF
C533 pgxor2 A_2 0.11fF
C534 S1 gnd 0.07fF
C535 S0 gnd 0.89fF
C536 a_156_n58# S0 0.17fF
C537 w_38_n97# C0bar 0.21fF
C538 G3 w_38_n424# 0.06fF
C539 a_44_n440# gnd 0.12fF
C540 GPG1 P32 0.09fF
C541 P10 GPG3 0.05fF
C542 pgxor2 a_n101_n282# 0.12fF
C543 a_254_n252# w_137_n280# 0.11fF
C544 Gout gnd 0.03fF
C545 clk a_278_n59# 0.33fF
C546 clk w_137_n171# 0.37fF
C547 a_254_n59# gnd 0.08fF
C548 a_75_n440# VDD 0.08fF
C549 a_75_n222# w_38_n206# 0.10fF
C550 C2 VDD 0.09fF
C551 a_296_n378# VDD 0.01fF
C552 w_137_n171# VDD 0.42fF
C553 a_333_n98# w_243_n62# 0.02fF
C554 a_278_n59# VDD 0.08fF
C555 s_0 C1 0.26fF
C556 a_318_n160# VDD 0.01fF
C557 a_84_n59# C0 0.16fF
C558 Pout w_38_n424# 0.05fF
C559 w_243_n62# a_300_n79# 0.09fF
C560 A_1 Pt1 0.09fF
C561 a_150_n274# w_137_n280# 0.15fF
C562 S3 a_149_n229# 0.04fF
C563 G3 w_n131_n463# 0.06fF
C564 a_150_n165# w_137_n171# 0.15fF
C565 pgxor2 w_n47_n271# 0.07fF
C566 a_150_n274# C1 0.04fF
C567 GPG1 pgxor2 0.05fF
C568 a_195_n452# VDD 0.02fF
C569 a_51_n200# VDD 0.01fF
C570 A_1 w_n47_n162# 0.19fF
C571 P21 GPG2 0.17fF
C572 S3 a_296_n269# 0.01fF
C573 a_150_n274# a_174_n296# 0.04fF
C574 C4 a_216_n386# 0.17fF
C575 P10 Pout 0.02fF
C576 S3 clk 0.19fF
C577 a_91_n232# gnd 0.02fF
C578 GPG1 G1 0.06fF
C579 Pt2 pgxor3 0.27fF
C580 w_143_n351# VDD 0.02fF
C581 B_2 gnd 0.11fF
C582 gnd a_44_n123# 0.11fF
C583 S3 VDD 1.07fF
C584 A_0 C0bar 0.10fF
C585 GPG2 w_38_n315# 0.19fF
C586 Pt2 w_38_n424# 0.14fF
C587 w_38_n97# Pt0 0.12fF
C588 C3 gnd 0.02fF
C589 G3 a_n30_n423# 0.02fF
C590 A_2 VDD 0.28fF
C591 clk w_243_n364# 0.37fF
C592 VDD a_75_n113# 0.02fF
C593 C0 a_44_n123# 0.07fF
C594 Pt2 G2 0.85fF
C595 w_243_n364# VDD 0.12fF
C596 a_156_n58# gnd 0.08fF
C597 P10 P21 0.04fF
C598 P10 w_38_n206# 0.07fF
C599 C0 gnd 0.33fF
C600 G2 w_38_n315# 0.06fF
C601 C1 w_123_n108# 0.40fF
C602 s_2 gnd 0.02fF
C603 w_38_n97# VDD 0.27fF
C604 a_44_n331# a_75_n331# 0.04fF
C605 GPG1 w_137_n389# 0.12fF
C606 pgxor2 G1 0.75fF
C607 a_174_n187# gnd 0.02fF
C608 Pt0 C0bar 0.07fF
C609 s_1 S1 0.06fF
C610 a_189_n117# VDD 0.01fF
C611 clk a_180_n58# 0.33fF
C612 pgxor1 S0 0.03fF
C613 s_1 S0 0.11fF
C614 GPG1 VDD 0.14fF
C615 Cout gnd 0.15fF
C616 G2 w_n131_n354# 0.06fF
C617 P32 w_137_n389# 0.06fF
C618 a_180_n58# VDD 0.08fF
C619 A_3 gnd 0.07fF
C620 w_243_n62# a_278_n59# 0.12fF
C621 B_1 A_1 0.32fF
C622 A_0 Pt0 0.09fF
C623 a_n101_n391# gnd 0.28fF
C624 a_150_n165# GPG1 0.07fF
C625 P32 VDD 0.32fF
C626 Pt1 P21 0.28fF
C627 a_136_n124# gnd 0.42fF
C628 a_183_n187# C2 0.04fF
C629 Pt1 w_38_n206# 0.25fF
C630 a_183_n187# w_137_n171# 0.10fF
C631 Pt1 Pt2 0.07fF
C632 a_44_n440# w_38_n424# 0.10fF
C633 C0bar VDD 1.23fF
C634 a_296_n76# VDD 0.01fF
C635 a_216_n386# w_189_n473# 0.03fF
C636 a_150_n415# gnd 0.02fF
C637 Pt1 w_n131_n245# 0.04fF
C638 G0 a_75_n113# 0.09fF
C639 Pt1 w_38_n315# 0.14fF
C640 a_278_n252# S3 0.12fF
C641 Pout Gnd 0.45fF
C642 a_195_n452# Gnd 0.16fF
C643 a_216_n386# Gnd 0.19fF
C644 Gout Gnd 0.14fF
C645 G3 Gnd 0.43fF
C646 a_75_n440# Gnd 0.13fF
C647 a_44_n440# Gnd 0.02fF
C648 a_n101_n391# Gnd 0.26fF
C649 Pt3 Gnd 1.11fF
C650 GPG3 Gnd 0.92fF
C651 a_174_n405# Gnd 0.09fF
C652 a_150_n383# Gnd 0.09fF
C653 P32 Gnd 0.60fF
C654 A_3 Gnd 0.43fF
C655 B_3 Gnd 0.74fF
C656 C4 Gnd 0.04fF
C657 a_300_n381# Gnd 0.16fF
C658 a_278_n361# Gnd 0.13fF
C659 a_254_n361# Gnd 0.15fF
C660 G2 Gnd 0.99fF
C661 a_75_n331# Gnd 0.13fF
C662 a_44_n331# Gnd 0.06fF
C663 a_n101_n282# Gnd 0.26fF
C664 pgxor3 Gnd 2.60fF
C665 a_231_n296# Gnd 0.21fF
C666 Pt2 Gnd 1.65fF
C667 C3 Gnd 0.02fF
C668 a_183_n296# Gnd 0.13fF
C669 GPG2 Gnd 0.57fF
C670 a_174_n296# Gnd 0.09fF
C671 a_150_n274# Gnd 0.09fF
C672 P21 Gnd 0.05fF
C673 A_2 Gnd 0.43fF
C674 B_2 Gnd 0.74fF
C675 a_149_n229# Gnd 0.02fF
C676 s_3 Gnd 0.18fF
C677 a_300_n272# Gnd 0.16fF
C678 S3 Gnd 0.00fF
C679 a_278_n252# Gnd 0.13fF
C680 a_254_n252# Gnd 0.15fF
C681 G1 Gnd 0.98fF
C682 a_75_n222# Gnd 0.13fF
C683 a_44_n222# Gnd 0.06fF
C684 a_n101_n173# Gnd 0.26fF
C685 pgxor2 Gnd 2.56fF
C686 Pt1 Gnd 1.65fF
C687 a_183_n187# Gnd 0.15fF
C688 GPG1 Gnd 1.38fF
C689 a_174_n187# Gnd 0.09fF
C690 a_150_n165# Gnd 0.09fF
C691 P10 Gnd 0.04fF
C692 A_1 Gnd 0.43fF
C693 B_1 Gnd 0.74fF
C694 a_153_n133# Gnd 0.02fF
C695 a_189_n117# Gnd 0.02fF
C696 s_2 Gnd 0.18fF
C697 a_300_n163# Gnd 0.16fF
C698 S2 Gnd 0.27fF
C699 a_278_n143# Gnd 0.13fF
C700 a_254_n143# Gnd 0.12fF
C701 a_333_n98# Gnd 0.02fF
C702 a_136_n124# Gnd 0.04fF
C703 pgxor1 Gnd 1.15fF
C704 C1 Gnd 0.55fF
C705 a_75_n113# Gnd 0.13fF
C706 G0 Gnd 0.00fF
C707 a_n101_n64# Gnd 0.26fF
C708 Pt0 Gnd 1.37fF
C709 s_1 Gnd 0.78fF
C710 a_300_n79# Gnd 0.16fF
C711 S1 Gnd 0.03fF
C712 s_0 Gnd 0.38fF
C713 a_202_n78# Gnd 0.16fF
C714 a_278_n59# Gnd 0.13fF
C715 a_254_n59# Gnd 0.15fF
C716 gnd Gnd 10.91fF
C717 S0 Gnd 0.03fF
C718 a_84_n59# Gnd 0.21fF
C719 A_0 Gnd 0.42fF
C720 B_0 Gnd 0.74fF
C721 C0bar Gnd 8.27fF
C722 C0 Gnd 2.30fF
C723 VDD Gnd 0.01fF
C724 pgxor0 Gnd 0.43fF
C725 a_180_n58# Gnd 0.13fF
C726 a_156_n58# Gnd 0.12fF
C727 clk Gnd 0.10fF
C728 w_189_n473# Gnd 2.44fF
C729 w_243_n364# Gnd 4.00fF
C730 w_137_n389# Gnd 4.21fF
C731 w_38_n424# Gnd 0.74fF
C732 w_n131_n463# Gnd 5.27fF
C733 w_n47_n380# Gnd 0.82fF
C734 w_143_n351# Gnd 0.17fF
C735 w_38_n315# Gnd 0.96fF
C736 w_n131_n354# Gnd 5.27fF
C737 w_n47_n271# Gnd 0.82fF
C738 w_137_n280# Gnd 0.04fF
C739 w_143_n242# Gnd 0.14fF
C740 w_205_n123# Gnd 0.77fF
C741 w_137_n171# Gnd 0.43fF
C742 w_38_n206# Gnd 0.69fF
C743 w_n131_n245# Gnd 5.27fF
C744 w_n47_n162# Gnd 0.82fF
C745 w_243_n62# Gnd 0.80fF
C746 w_123_n108# Gnd 0.31fF
C747 w_n47_n53# Gnd 0.82fF
C748 w_n131_n136# Gnd 6.10fF
C749 w_38_n97# Gnd 4.57fF


.tran 1n 100n
* .ic V(A_0) =0
* .ic V(A_1) =0
* .ic V(A_2) =0
* .ic V(A_3) =0

* .ic V(B_0) =0
* .ic V(B_1) =0
* .ic V(B_2) =0
* .ic V(B_3) =0

* .ic V(C0) =0

.ic V(S0)=0
.ic V(S1)=0
.ic V(S2)=0
.ic V(S3)=0

.ic V(Cout) =0


* 'SUPPLY'

* V1 A0 gnd 'SUPPLY'
* V2 A1 gnd 0
* V3 A2 gnd 0
* V4 A3 gnd 0

* V5 B0 gnd 0
* V6 B1 gnd 0
* V7 B2 gnd 0
* V8 B3 gnd 0

* V9 C0 gnd 0

V1 A_0 gnd 0    
* V1 A_0 gnd 'SUPPLY'
V2 A_1 gnd 0
* V2 A_1 gnd 'SUPPLY'
V3 A_2 gnd 0
* V3 A_2 gnd 'SUPPLY'
V4 A_3 gnd 0
* V4 A_3 gnd 'SUPPLY'

* V5 B_0 gnd 0
V5 B_0 gnd 'SUPPLY'
V6 B_1 gnd 0
* V6 B_1 gnd 'SUPPLY'
V7 B_2 gnd 0
* V7 B_2 gnd 'SUPPLY'
V8 B_3 gnd 0
* V8 B_3 gnd 'SUPPLY'
* * V5 B_0 gnd PULSE(0 'SUPPLY' 50ns 50ps 50ps 30ns 60ns)
* V1 A0 gnd PULSE(0 'SUPPLY' 20ns 10ps 10ps 30ns 60ns)
V10 clk gnd PULSE(0 'SUPPLY' 30ns 10ps 10ps 30ns 60ns)

V9 C0 gnd 0
* V9 C0 gnd 'SUPPLY'
* * V10 clk gnd 'SUPPLY'

* .measure tran B0_val FIND v(B_0) AT=8n
* .measure tran S0_val FIND v(s_0) AT=8n
* .measure tran S1_val FIND v(s_1) AT=8n
* .measure tran S2_val FIND v(s_2) AT=8n  
* .measure tran S3_val FIND v(s_3) AT=8n  
* .measure tran C4_val FIND v(C4) AT=8n
* .measure tran C0_val FIND v(C0) AT=8n
* .measure tran C2_val FIND v(C2) AT=8n
* .measure tran C3_val FIND v(C3) AT=8n
* .measure tran G0_val FIND v(G0) AT=8n
* .measure tran G2_val FIND v(G2) AT=8n
* .measure tran P2_val FIND v(Pt2) AT=8n
* .measure tran P21 FIND v(P21) AT=8n
* .measure tran P10 FIND v(P10) AT=8n
* .measure tran P1_val FIND v(Pt1) AT=8n
* .measure tran GPG2_val FIND v(GPG2) AT=8n
 
.control
run
plot V(s_0)+6 V(S0)+3 V(S1) V(clk)-3
.endc