magic
tech scmos
timestamp 1731351332
<< nwell >>
rect -21 8 31 60
<< ntransistor >>
rect -10 -9 -8 2
rect 12 -9 14 2
<< ptransistor >>
rect -10 14 -8 54
rect -4 14 -2 54
rect 12 14 14 54
rect 18 14 20 54
<< ndiffusion >>
rect -15 -5 -10 2
rect -11 -9 -10 -5
rect -8 -2 -7 2
rect -8 -9 -3 -2
rect 7 -5 12 2
rect 11 -9 12 -5
rect 14 -2 15 2
rect 14 -9 19 -2
<< pdiffusion >>
rect -11 50 -10 54
rect -15 14 -10 50
rect -8 14 -4 54
rect -2 18 3 54
rect -2 14 -1 18
rect 11 50 12 54
rect 7 14 12 50
rect 14 14 18 54
rect 20 18 25 54
rect 20 14 21 18
<< ndcontact >>
rect -15 -9 -11 -5
rect -7 -2 -3 2
rect 7 -9 11 -5
rect 15 -2 19 2
<< pdcontact >>
rect -15 50 -11 54
rect -1 14 3 18
rect 7 50 11 54
rect 21 14 25 18
<< polysilicon >>
rect -10 54 -8 57
rect -4 54 -2 65
rect 12 54 14 57
rect 18 54 20 65
rect -10 2 -8 14
rect -4 11 -2 14
rect 12 2 14 14
rect 18 11 20 14
rect -10 -12 -8 -9
rect 12 -12 14 -9
<< polycontact >>
rect -2 61 2 65
rect 14 61 18 65
rect -14 3 -10 7
rect 8 3 12 7
<< metal1 >>
rect 2 62 14 65
rect -14 55 10 58
rect -14 54 -11 55
rect 7 54 10 55
rect 0 7 3 14
rect 22 7 25 14
rect -20 4 -14 7
rect 0 4 8 7
rect 0 2 3 4
rect 22 4 31 7
rect 22 2 25 4
rect -3 -1 3 2
rect 19 -1 25 2
rect -15 -12 -12 -9
rect 7 -12 10 -9
rect -15 -15 10 -12
<< labels >>
rlabel metal1 -19 5 -19 5 3 D
rlabel metal1 -13 56 -13 56 1 VDD
rlabel metal1 7 63 7 63 5 clk
rlabel metal1 1 -14 1 -14 1 gnd
rlabel metal1 29 6 29 6 7 out
<< end >>
