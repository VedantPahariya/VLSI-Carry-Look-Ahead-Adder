magic
tech scmos
timestamp 1731492129
<< nwell >>
rect -152 -77 -64 -45
<< ntransistor >>
rect -141 -103 -139 -83
rect -133 -103 -131 -83
rect -117 -93 -115 -83
rect -101 -93 -99 -83
rect -93 -93 -91 -83
rect -77 -93 -75 -83
<< ptransistor >>
rect -141 -71 -139 -51
rect -133 -71 -131 -51
rect -117 -71 -115 -51
rect -101 -71 -99 -51
rect -93 -71 -91 -51
rect -77 -71 -75 -51
<< ndiffusion >>
rect -146 -99 -141 -83
rect -142 -103 -141 -99
rect -139 -103 -133 -83
rect -131 -87 -130 -83
rect -131 -103 -126 -87
rect -122 -89 -117 -83
rect -118 -93 -117 -89
rect -115 -87 -114 -83
rect -115 -93 -110 -87
rect -102 -87 -101 -83
rect -106 -93 -101 -87
rect -99 -89 -93 -83
rect -99 -93 -98 -89
rect -94 -93 -93 -89
rect -91 -87 -90 -83
rect -91 -93 -86 -87
rect -82 -89 -77 -83
rect -78 -93 -77 -89
rect -75 -87 -74 -83
rect -75 -93 -70 -87
<< pdiffusion >>
rect -142 -55 -141 -51
rect -146 -71 -141 -55
rect -139 -67 -133 -51
rect -139 -71 -138 -67
rect -134 -71 -133 -67
rect -131 -55 -130 -51
rect -131 -71 -126 -55
rect -118 -55 -117 -51
rect -122 -71 -117 -55
rect -115 -67 -110 -51
rect -115 -71 -114 -67
rect -102 -55 -101 -51
rect -106 -71 -101 -55
rect -99 -71 -93 -51
rect -91 -67 -86 -51
rect -91 -71 -90 -67
rect -78 -55 -77 -51
rect -82 -71 -77 -55
rect -75 -67 -70 -51
rect -75 -71 -74 -67
<< ndcontact >>
rect -146 -103 -142 -99
rect -130 -87 -126 -83
rect -122 -93 -118 -89
rect -114 -87 -110 -83
rect -106 -87 -102 -83
rect -98 -93 -94 -89
rect -90 -87 -86 -83
rect -82 -93 -78 -89
rect -74 -87 -70 -83
<< pdcontact >>
rect -146 -55 -142 -51
rect -138 -71 -134 -67
rect -130 -55 -126 -51
rect -122 -55 -118 -51
rect -114 -71 -110 -67
rect -106 -55 -102 -51
rect -90 -71 -86 -67
rect -82 -55 -78 -51
rect -74 -71 -70 -67
<< polysilicon >>
rect -141 -51 -139 -48
rect -133 -51 -131 -48
rect -117 -51 -115 -48
rect -101 -51 -99 -48
rect -93 -51 -91 -48
rect -77 -51 -75 -48
rect -141 -83 -139 -71
rect -133 -83 -131 -71
rect -117 -83 -115 -71
rect -101 -83 -99 -71
rect -93 -75 -91 -71
rect -93 -83 -91 -80
rect -77 -83 -75 -71
rect -117 -96 -115 -93
rect -101 -96 -99 -93
rect -93 -96 -91 -93
rect -77 -96 -75 -93
rect -141 -106 -139 -103
rect -133 -105 -131 -103
<< polycontact >>
rect -145 -76 -141 -72
rect -121 -76 -117 -72
rect -105 -76 -101 -72
rect -81 -82 -77 -78
rect -135 -109 -131 -105
<< metal1 >>
rect -152 -48 -64 -45
rect -146 -51 -143 -48
rect -129 -51 -126 -48
rect -122 -51 -119 -48
rect -106 -51 -103 -48
rect -82 -51 -79 -48
rect -86 -71 -82 -68
rect -159 -76 -145 -73
rect -137 -73 -134 -71
rect -137 -76 -121 -73
rect -113 -73 -110 -71
rect -113 -76 -105 -73
rect -129 -83 -126 -76
rect -113 -83 -110 -76
rect -85 -78 -82 -71
rect -73 -78 -70 -71
rect -85 -82 -81 -78
rect -73 -81 -58 -78
rect -85 -83 -82 -82
rect -73 -83 -70 -81
rect -102 -86 -90 -83
rect -86 -86 -82 -83
rect -122 -96 -119 -93
rect -97 -96 -94 -93
rect -82 -96 -79 -93
rect -146 -99 -79 -96
rect -158 -109 -135 -106
<< pm12contact >>
rect -93 -80 -88 -75
<< metal2 >>
rect -159 -80 -93 -77
<< labels >>
rlabel metal1 -140 -46 -140 -46 5 VDD
rlabel metal1 -102 -98 -102 -98 1 gnd
rlabel metal1 -72 -80 -72 -80 1 out
rlabel metal1 -158 -75 -158 -75 1 lastandC
rlabel metal1 -157 -108 -157 -108 1 lastandnr
rlabel metal2 -158 -79 -158 -79 1 lastORnd
<< end >>
