magic
tech scmos
timestamp 1731529929
<< nwell >>
rect 95 -7 136 -4
rect 71 -24 136 -7
rect -131 -51 -107 -31
rect -131 -63 -75 -51
rect -47 -53 -6 -33
rect 71 -39 95 -24
rect -107 -77 -75 -63
rect 38 -65 71 -45
rect -94 -92 -36 -77
rect -94 -104 -39 -92
rect 38 -97 110 -65
rect 143 -76 188 -73
rect 123 -93 188 -76
rect -131 -136 -39 -104
rect 123 -108 147 -93
rect -47 -162 -6 -142
rect -107 -186 -75 -162
rect 70 -174 102 -137
rect 131 -171 219 -139
rect 249 -142 290 -139
rect 225 -159 290 -142
rect 225 -174 249 -159
rect -94 -201 -36 -186
rect -94 -213 -39 -201
rect 38 -206 110 -174
rect -131 -245 -39 -213
rect -47 -271 -6 -251
rect -107 -295 -75 -271
rect 70 -283 102 -246
rect 131 -280 219 -248
rect 249 -251 290 -248
rect 225 -268 290 -251
rect 225 -283 249 -268
rect -94 -310 -36 -295
rect -94 -322 -39 -310
rect 38 -315 110 -283
rect -131 -354 -39 -322
rect -47 -380 -6 -360
rect -107 -404 -75 -380
rect -94 -419 -36 -404
rect -94 -431 -39 -419
rect 38 -424 110 -392
rect -131 -463 -39 -431
<< ntransistor >>
rect 106 -34 108 -30
rect 122 -34 124 -30
rect -36 -63 -34 -59
rect -20 -63 -18 -59
rect -69 -66 -59 -64
rect -120 -79 -118 -69
rect -30 -90 10 -88
rect 82 -55 84 -45
rect -30 -98 10 -96
rect -33 -117 7 -115
rect 49 -123 51 -103
rect 57 -123 59 -103
rect 73 -113 75 -103
rect 89 -123 91 -103
rect 97 -123 99 -103
rect 158 -103 160 -99
rect 174 -103 176 -99
rect -33 -125 7 -123
rect 134 -124 136 -114
rect 54 -150 64 -148
rect 54 -158 64 -156
rect -36 -172 -34 -168
rect -20 -172 -18 -168
rect -69 -175 -59 -173
rect -30 -199 10 -197
rect 142 -197 144 -177
rect 150 -197 152 -177
rect 166 -187 168 -177
rect 182 -187 184 -177
rect 190 -187 192 -177
rect 206 -187 208 -177
rect 260 -169 262 -165
rect 276 -169 278 -165
rect 236 -190 238 -180
rect -30 -207 10 -205
rect 49 -222 51 -212
rect 57 -222 59 -212
rect 73 -222 75 -212
rect -33 -226 7 -224
rect 89 -232 91 -212
rect 97 -232 99 -212
rect -33 -234 7 -232
rect 54 -259 64 -257
rect 54 -267 64 -265
rect -36 -281 -34 -277
rect -20 -281 -18 -277
rect -69 -284 -59 -282
rect -30 -308 10 -306
rect 142 -306 144 -286
rect 150 -306 152 -286
rect 166 -296 168 -286
rect 182 -296 184 -286
rect 190 -296 192 -286
rect 206 -296 208 -286
rect 260 -278 262 -274
rect 276 -278 278 -274
rect 236 -299 238 -289
rect -30 -316 10 -314
rect 49 -331 51 -321
rect 57 -331 59 -321
rect 73 -331 75 -321
rect -33 -335 7 -333
rect 89 -341 91 -321
rect 97 -341 99 -321
rect -33 -343 7 -341
rect -36 -390 -34 -386
rect -20 -390 -18 -386
rect -69 -393 -59 -391
rect -30 -417 10 -415
rect -30 -425 10 -423
rect 49 -440 51 -430
rect 57 -440 59 -430
rect 73 -440 75 -430
rect -33 -444 7 -442
rect 89 -450 91 -430
rect 97 -450 99 -430
rect -33 -452 7 -450
<< ptransistor >>
rect 82 -33 84 -13
rect 106 -18 108 -10
rect 122 -18 124 -10
rect -120 -57 -118 -37
rect -36 -47 -34 -39
rect -20 -47 -18 -39
rect -101 -66 -81 -64
rect -88 -90 -48 -88
rect 49 -91 51 -51
rect 57 -91 59 -51
rect 73 -91 75 -71
rect 89 -91 91 -71
rect 97 -91 99 -71
rect -88 -98 -48 -96
rect 134 -102 136 -82
rect 158 -87 160 -79
rect 174 -87 176 -79
rect -125 -117 -45 -115
rect -125 -125 -45 -123
rect -36 -156 -34 -148
rect -20 -156 -18 -148
rect 76 -150 96 -148
rect 76 -158 96 -156
rect 142 -165 144 -145
rect 150 -165 152 -145
rect 166 -165 168 -145
rect 182 -165 184 -145
rect 190 -165 192 -145
rect 206 -165 208 -145
rect -101 -175 -81 -173
rect 236 -168 238 -148
rect 260 -153 262 -145
rect 276 -153 278 -145
rect -88 -199 -48 -197
rect 49 -200 51 -180
rect 57 -200 59 -180
rect 73 -200 75 -180
rect 89 -200 91 -180
rect 97 -200 99 -180
rect -88 -207 -48 -205
rect -125 -226 -45 -224
rect -125 -234 -45 -232
rect -36 -265 -34 -257
rect -20 -265 -18 -257
rect 76 -259 96 -257
rect 76 -267 96 -265
rect 142 -274 144 -254
rect 150 -274 152 -254
rect 166 -274 168 -254
rect 182 -274 184 -254
rect 190 -274 192 -254
rect 206 -274 208 -254
rect -101 -284 -81 -282
rect 236 -277 238 -257
rect 260 -262 262 -254
rect 276 -262 278 -254
rect -88 -308 -48 -306
rect 49 -309 51 -289
rect 57 -309 59 -289
rect 73 -309 75 -289
rect 89 -309 91 -289
rect 97 -309 99 -289
rect -88 -316 -48 -314
rect -125 -335 -45 -333
rect -125 -343 -45 -341
rect -36 -374 -34 -366
rect -20 -374 -18 -366
rect -101 -393 -81 -391
rect -88 -417 -48 -415
rect 49 -418 51 -398
rect 57 -418 59 -398
rect 73 -418 75 -398
rect 89 -418 91 -398
rect 97 -418 99 -398
rect -88 -425 -48 -423
rect -125 -444 -45 -442
rect -125 -452 -45 -450
<< ndiffusion >>
rect 105 -34 106 -30
rect 108 -34 109 -30
rect 121 -34 122 -30
rect 124 -34 125 -30
rect 77 -51 82 -45
rect -65 -63 -59 -59
rect -37 -63 -36 -59
rect -34 -63 -33 -59
rect -21 -63 -20 -59
rect -18 -63 -17 -59
rect -69 -64 -59 -63
rect -125 -75 -120 -69
rect -121 -79 -120 -75
rect -118 -73 -117 -69
rect -69 -67 -59 -66
rect -69 -71 -63 -67
rect -118 -79 -113 -73
rect -26 -87 10 -83
rect -30 -88 10 -87
rect -30 -96 10 -90
rect 81 -55 82 -51
rect 84 -49 85 -45
rect 84 -55 89 -49
rect -30 -99 10 -98
rect -30 -103 6 -99
rect 48 -107 49 -103
rect -29 -114 7 -110
rect -33 -115 7 -114
rect -33 -118 7 -117
rect -33 -122 3 -118
rect -33 -123 7 -122
rect 44 -123 49 -107
rect 51 -119 57 -103
rect 51 -123 52 -119
rect 56 -123 57 -119
rect 59 -107 60 -103
rect 59 -123 64 -107
rect 68 -109 73 -103
rect 72 -113 73 -109
rect 75 -107 76 -103
rect 75 -113 80 -107
rect 84 -119 89 -103
rect 88 -123 89 -119
rect 91 -123 97 -103
rect 99 -107 100 -103
rect 99 -123 104 -107
rect 157 -103 158 -99
rect 160 -103 161 -99
rect 173 -103 174 -99
rect 176 -103 177 -99
rect 129 -120 134 -114
rect -33 -126 7 -125
rect 133 -124 134 -120
rect 136 -118 137 -114
rect 136 -124 141 -118
rect -29 -130 7 -126
rect 54 -147 60 -143
rect 54 -148 64 -147
rect 54 -151 64 -150
rect 58 -155 64 -151
rect 54 -156 64 -155
rect 54 -159 64 -158
rect 54 -163 60 -159
rect -65 -172 -59 -168
rect -37 -172 -36 -168
rect -34 -172 -33 -168
rect -21 -172 -20 -168
rect -18 -172 -17 -168
rect -69 -173 -59 -172
rect -69 -176 -59 -175
rect -69 -180 -63 -176
rect -26 -196 10 -192
rect -30 -197 10 -196
rect -30 -205 10 -199
rect 137 -193 142 -177
rect 141 -197 142 -193
rect 144 -197 150 -177
rect 152 -181 153 -177
rect 152 -197 157 -181
rect 161 -183 166 -177
rect 165 -187 166 -183
rect 168 -181 169 -177
rect 168 -187 173 -181
rect 181 -181 182 -177
rect 177 -187 182 -181
rect 184 -183 190 -177
rect 184 -187 185 -183
rect 189 -187 190 -183
rect 192 -181 193 -177
rect 192 -187 197 -181
rect 201 -183 206 -177
rect 205 -187 206 -183
rect 208 -181 209 -177
rect 259 -169 260 -165
rect 262 -169 263 -165
rect 275 -169 276 -165
rect 278 -169 279 -165
rect 208 -187 213 -181
rect 231 -186 236 -180
rect 235 -190 236 -186
rect 238 -184 239 -180
rect 238 -190 243 -184
rect -30 -208 10 -207
rect -30 -212 6 -208
rect 48 -216 49 -212
rect -29 -223 7 -219
rect 44 -222 49 -216
rect 51 -218 57 -212
rect 51 -222 52 -218
rect 56 -222 57 -218
rect 59 -216 60 -212
rect 59 -222 64 -216
rect 68 -218 73 -212
rect 72 -222 73 -218
rect 75 -216 76 -212
rect 75 -222 80 -216
rect -33 -224 7 -223
rect -33 -227 7 -226
rect -33 -231 3 -227
rect -33 -232 7 -231
rect 84 -228 89 -212
rect 88 -232 89 -228
rect 91 -232 97 -212
rect 99 -216 100 -212
rect 99 -232 104 -216
rect -33 -235 7 -234
rect -29 -239 7 -235
rect 54 -256 60 -252
rect 54 -257 64 -256
rect 54 -260 64 -259
rect 58 -264 64 -260
rect 54 -265 64 -264
rect 54 -268 64 -267
rect 54 -272 60 -268
rect -65 -281 -59 -277
rect -37 -281 -36 -277
rect -34 -281 -33 -277
rect -21 -281 -20 -277
rect -18 -281 -17 -277
rect -69 -282 -59 -281
rect -69 -285 -59 -284
rect -69 -289 -63 -285
rect -26 -305 10 -301
rect -30 -306 10 -305
rect -30 -314 10 -308
rect 137 -302 142 -286
rect 141 -306 142 -302
rect 144 -306 150 -286
rect 152 -290 153 -286
rect 152 -306 157 -290
rect 161 -292 166 -286
rect 165 -296 166 -292
rect 168 -290 169 -286
rect 168 -296 173 -290
rect 181 -290 182 -286
rect 177 -296 182 -290
rect 184 -292 190 -286
rect 184 -296 185 -292
rect 189 -296 190 -292
rect 192 -290 193 -286
rect 192 -296 197 -290
rect 201 -292 206 -286
rect 205 -296 206 -292
rect 208 -290 209 -286
rect 259 -278 260 -274
rect 262 -278 263 -274
rect 275 -278 276 -274
rect 278 -278 279 -274
rect 208 -296 213 -290
rect 231 -295 236 -289
rect 235 -299 236 -295
rect 238 -293 239 -289
rect 238 -299 243 -293
rect -30 -317 10 -316
rect -30 -321 6 -317
rect 48 -325 49 -321
rect -29 -332 7 -328
rect 44 -331 49 -325
rect 51 -327 57 -321
rect 51 -331 52 -327
rect 56 -331 57 -327
rect 59 -325 60 -321
rect 59 -331 64 -325
rect 68 -327 73 -321
rect 72 -331 73 -327
rect 75 -325 76 -321
rect 75 -331 80 -325
rect -33 -333 7 -332
rect -33 -336 7 -335
rect -33 -340 3 -336
rect -33 -341 7 -340
rect 84 -337 89 -321
rect 88 -341 89 -337
rect 91 -341 97 -321
rect 99 -325 100 -321
rect 99 -341 104 -325
rect -33 -344 7 -343
rect -29 -348 7 -344
rect -65 -390 -59 -386
rect -37 -390 -36 -386
rect -34 -390 -33 -386
rect -21 -390 -20 -386
rect -18 -390 -17 -386
rect -69 -391 -59 -390
rect -69 -394 -59 -393
rect -69 -398 -63 -394
rect -26 -414 10 -410
rect -30 -415 10 -414
rect -30 -423 10 -417
rect -30 -426 10 -425
rect -30 -430 6 -426
rect 48 -434 49 -430
rect -29 -441 7 -437
rect 44 -440 49 -434
rect 51 -436 57 -430
rect 51 -440 52 -436
rect 56 -440 57 -436
rect 59 -434 60 -430
rect 59 -440 64 -434
rect 68 -436 73 -430
rect 72 -440 73 -436
rect 75 -434 76 -430
rect 75 -440 80 -434
rect -33 -442 7 -441
rect -33 -445 7 -444
rect -33 -449 3 -445
rect -33 -450 7 -449
rect 84 -446 89 -430
rect 88 -450 89 -446
rect 91 -450 97 -430
rect 99 -434 100 -430
rect 99 -450 104 -434
rect -33 -453 7 -452
rect -29 -457 7 -453
<< pdiffusion >>
rect 81 -17 82 -13
rect 77 -33 82 -17
rect 84 -29 89 -13
rect 101 -14 106 -10
rect 105 -18 106 -14
rect 108 -14 113 -10
rect 108 -18 109 -14
rect 117 -14 122 -10
rect 121 -18 122 -14
rect 124 -13 129 -10
rect 124 -18 125 -13
rect 84 -33 85 -29
rect -121 -41 -120 -37
rect -125 -57 -120 -41
rect -118 -53 -113 -37
rect -41 -43 -36 -39
rect -37 -47 -36 -43
rect -34 -43 -29 -39
rect -34 -47 -33 -43
rect -25 -43 -20 -39
rect -21 -47 -20 -43
rect -18 -42 -13 -39
rect -18 -47 -17 -42
rect -118 -57 -117 -53
rect 48 -55 49 -51
rect -101 -63 -85 -59
rect -101 -64 -81 -63
rect -101 -67 -81 -66
rect -97 -71 -81 -67
rect -84 -87 -48 -83
rect -88 -88 -48 -87
rect -88 -91 -48 -90
rect -88 -95 -52 -91
rect -88 -96 -48 -95
rect 44 -91 49 -55
rect 51 -91 57 -51
rect 59 -87 64 -51
rect 59 -91 60 -87
rect 72 -75 73 -71
rect 68 -91 73 -75
rect 75 -87 80 -71
rect 75 -91 76 -87
rect 88 -75 89 -71
rect 84 -91 89 -75
rect 91 -87 97 -71
rect 91 -91 92 -87
rect 96 -91 97 -87
rect 99 -75 100 -71
rect 99 -91 104 -75
rect 133 -86 134 -82
rect -88 -99 -48 -98
rect -84 -103 -48 -99
rect 129 -102 134 -86
rect 136 -98 141 -82
rect 153 -83 158 -79
rect 157 -87 158 -83
rect 160 -83 165 -79
rect 160 -87 161 -83
rect 169 -83 174 -79
rect 173 -87 174 -83
rect 176 -82 181 -79
rect 176 -87 177 -82
rect 136 -102 137 -98
rect -121 -114 -45 -110
rect -125 -115 -45 -114
rect -125 -123 -45 -117
rect -125 -126 -45 -125
rect -125 -130 -49 -126
rect -41 -152 -36 -148
rect -37 -156 -36 -152
rect -34 -152 -29 -148
rect -34 -156 -33 -152
rect -25 -152 -20 -148
rect -21 -156 -20 -152
rect -18 -151 -13 -148
rect 80 -147 96 -143
rect 76 -148 96 -147
rect 141 -149 142 -145
rect -18 -156 -17 -151
rect 76 -156 96 -150
rect 76 -159 96 -158
rect 76 -163 92 -159
rect 137 -165 142 -149
rect 144 -161 150 -145
rect 144 -165 145 -161
rect 149 -165 150 -161
rect 152 -149 153 -145
rect 152 -165 157 -149
rect 165 -149 166 -145
rect 161 -165 166 -149
rect 168 -161 173 -145
rect 168 -165 169 -161
rect 181 -149 182 -145
rect 177 -165 182 -149
rect 184 -165 190 -145
rect 192 -161 197 -145
rect 192 -165 193 -161
rect 205 -149 206 -145
rect 201 -165 206 -149
rect 208 -161 213 -145
rect 208 -165 209 -161
rect 235 -152 236 -148
rect -101 -172 -85 -168
rect -101 -173 -81 -172
rect -101 -176 -81 -175
rect -97 -180 -81 -176
rect 231 -168 236 -152
rect 238 -164 243 -148
rect 255 -149 260 -145
rect 259 -153 260 -149
rect 262 -149 267 -145
rect 262 -153 263 -149
rect 271 -149 276 -145
rect 275 -153 276 -149
rect 278 -148 283 -145
rect 278 -153 279 -148
rect 238 -168 239 -164
rect 48 -184 49 -180
rect -84 -196 -48 -192
rect -88 -197 -48 -196
rect -88 -200 -48 -199
rect -88 -204 -52 -200
rect -88 -205 -48 -204
rect 44 -200 49 -184
rect 51 -200 57 -180
rect 59 -196 64 -180
rect 59 -200 60 -196
rect 72 -184 73 -180
rect 68 -200 73 -184
rect 75 -196 80 -180
rect 75 -200 76 -196
rect 88 -184 89 -180
rect 84 -200 89 -184
rect 91 -196 97 -180
rect 91 -200 92 -196
rect 96 -200 97 -196
rect 99 -184 100 -180
rect 99 -200 104 -184
rect -88 -208 -48 -207
rect -84 -212 -48 -208
rect -121 -223 -45 -219
rect -125 -224 -45 -223
rect -125 -232 -45 -226
rect -125 -235 -45 -234
rect -125 -239 -49 -235
rect -41 -261 -36 -257
rect -37 -265 -36 -261
rect -34 -261 -29 -257
rect -34 -265 -33 -261
rect -25 -261 -20 -257
rect -21 -265 -20 -261
rect -18 -260 -13 -257
rect 80 -256 96 -252
rect 76 -257 96 -256
rect 141 -258 142 -254
rect -18 -265 -17 -260
rect 76 -265 96 -259
rect 76 -268 96 -267
rect 76 -272 92 -268
rect 137 -274 142 -258
rect 144 -270 150 -254
rect 144 -274 145 -270
rect 149 -274 150 -270
rect 152 -258 153 -254
rect 152 -274 157 -258
rect 165 -258 166 -254
rect 161 -274 166 -258
rect 168 -270 173 -254
rect 168 -274 169 -270
rect 181 -258 182 -254
rect 177 -274 182 -258
rect 184 -274 190 -254
rect 192 -270 197 -254
rect 192 -274 193 -270
rect 205 -258 206 -254
rect 201 -274 206 -258
rect 208 -270 213 -254
rect 208 -274 209 -270
rect 235 -261 236 -257
rect -101 -281 -85 -277
rect -101 -282 -81 -281
rect -101 -285 -81 -284
rect -97 -289 -81 -285
rect 231 -277 236 -261
rect 238 -273 243 -257
rect 255 -258 260 -254
rect 259 -262 260 -258
rect 262 -258 267 -254
rect 262 -262 263 -258
rect 271 -258 276 -254
rect 275 -262 276 -258
rect 278 -257 283 -254
rect 278 -262 279 -257
rect 238 -277 239 -273
rect 48 -293 49 -289
rect -84 -305 -48 -301
rect -88 -306 -48 -305
rect -88 -309 -48 -308
rect -88 -313 -52 -309
rect -88 -314 -48 -313
rect 44 -309 49 -293
rect 51 -309 57 -289
rect 59 -305 64 -289
rect 59 -309 60 -305
rect 72 -293 73 -289
rect 68 -309 73 -293
rect 75 -305 80 -289
rect 75 -309 76 -305
rect 88 -293 89 -289
rect 84 -309 89 -293
rect 91 -305 97 -289
rect 91 -309 92 -305
rect 96 -309 97 -305
rect 99 -293 100 -289
rect 99 -309 104 -293
rect -88 -317 -48 -316
rect -84 -321 -48 -317
rect -121 -332 -45 -328
rect -125 -333 -45 -332
rect -125 -341 -45 -335
rect -125 -344 -45 -343
rect -125 -348 -49 -344
rect -41 -370 -36 -366
rect -37 -374 -36 -370
rect -34 -370 -29 -366
rect -34 -374 -33 -370
rect -25 -370 -20 -366
rect -21 -374 -20 -370
rect -18 -369 -13 -366
rect -18 -374 -17 -369
rect -101 -390 -85 -386
rect -101 -391 -81 -390
rect -101 -394 -81 -393
rect -97 -398 -81 -394
rect 48 -402 49 -398
rect -84 -414 -48 -410
rect -88 -415 -48 -414
rect -88 -418 -48 -417
rect -88 -422 -52 -418
rect -88 -423 -48 -422
rect 44 -418 49 -402
rect 51 -418 57 -398
rect 59 -414 64 -398
rect 59 -418 60 -414
rect 72 -402 73 -398
rect 68 -418 73 -402
rect 75 -414 80 -398
rect 75 -418 76 -414
rect 88 -402 89 -398
rect 84 -418 89 -402
rect 91 -414 97 -398
rect 91 -418 92 -414
rect 96 -418 97 -414
rect 99 -402 100 -398
rect 99 -418 104 -402
rect -88 -426 -48 -425
rect -84 -430 -48 -426
rect -121 -441 -45 -437
rect -125 -442 -45 -441
rect -125 -450 -45 -444
rect -125 -453 -45 -452
rect -125 -457 -49 -453
<< ndcontact >>
rect 101 -34 105 -30
rect 109 -34 113 -30
rect 117 -34 121 -30
rect -69 -63 -65 -59
rect -41 -63 -37 -59
rect -33 -63 -29 -59
rect -25 -63 -21 -59
rect -125 -79 -121 -75
rect -117 -73 -113 -69
rect -63 -71 -59 -67
rect -30 -87 -26 -83
rect 77 -55 81 -51
rect 85 -49 89 -45
rect 6 -103 10 -99
rect 44 -107 48 -103
rect -33 -114 -29 -110
rect 3 -122 7 -118
rect 52 -123 56 -119
rect 60 -107 64 -103
rect 68 -113 72 -109
rect 76 -107 80 -103
rect 84 -123 88 -119
rect 100 -107 104 -103
rect 153 -103 157 -99
rect 161 -103 165 -99
rect 169 -103 173 -99
rect 129 -124 133 -120
rect 137 -118 141 -114
rect -33 -130 -29 -126
rect 60 -147 64 -143
rect 54 -155 58 -151
rect 60 -163 64 -159
rect -69 -172 -65 -168
rect -41 -172 -37 -168
rect -33 -172 -29 -168
rect -25 -172 -21 -168
rect -63 -180 -59 -176
rect -30 -196 -26 -192
rect 137 -197 141 -193
rect 153 -181 157 -177
rect 161 -187 165 -183
rect 169 -181 173 -177
rect 177 -181 181 -177
rect 185 -187 189 -183
rect 193 -181 197 -177
rect 201 -187 205 -183
rect 209 -181 213 -177
rect 255 -169 259 -165
rect 263 -169 267 -165
rect 271 -169 275 -165
rect 231 -190 235 -186
rect 239 -184 243 -180
rect 6 -212 10 -208
rect 44 -216 48 -212
rect -33 -223 -29 -219
rect 52 -222 56 -218
rect 60 -216 64 -212
rect 68 -222 72 -218
rect 76 -216 80 -212
rect 3 -231 7 -227
rect 84 -232 88 -228
rect 100 -216 104 -212
rect -33 -239 -29 -235
rect 60 -256 64 -252
rect 54 -264 58 -260
rect 60 -272 64 -268
rect -69 -281 -65 -277
rect -41 -281 -37 -277
rect -33 -281 -29 -277
rect -25 -281 -21 -277
rect -63 -289 -59 -285
rect -30 -305 -26 -301
rect 137 -306 141 -302
rect 153 -290 157 -286
rect 161 -296 165 -292
rect 169 -290 173 -286
rect 177 -290 181 -286
rect 185 -296 189 -292
rect 193 -290 197 -286
rect 201 -296 205 -292
rect 209 -290 213 -286
rect 255 -278 259 -274
rect 263 -278 267 -274
rect 271 -278 275 -274
rect 231 -299 235 -295
rect 239 -293 243 -289
rect 6 -321 10 -317
rect 44 -325 48 -321
rect -33 -332 -29 -328
rect 52 -331 56 -327
rect 60 -325 64 -321
rect 68 -331 72 -327
rect 76 -325 80 -321
rect 3 -340 7 -336
rect 84 -341 88 -337
rect 100 -325 104 -321
rect -33 -348 -29 -344
rect -69 -390 -65 -386
rect -41 -390 -37 -386
rect -33 -390 -29 -386
rect -25 -390 -21 -386
rect -63 -398 -59 -394
rect -30 -414 -26 -410
rect 6 -430 10 -426
rect 44 -434 48 -430
rect -33 -441 -29 -437
rect 52 -440 56 -436
rect 60 -434 64 -430
rect 68 -440 72 -436
rect 76 -434 80 -430
rect 3 -449 7 -445
rect 84 -450 88 -446
rect 100 -434 104 -430
rect -33 -457 -29 -453
<< pdcontact >>
rect 77 -17 81 -13
rect 101 -18 105 -14
rect 109 -18 113 -14
rect 117 -18 121 -14
rect 85 -33 89 -29
rect -125 -41 -121 -37
rect -41 -47 -37 -43
rect -33 -47 -29 -43
rect -25 -47 -21 -43
rect -117 -57 -113 -53
rect 44 -55 48 -51
rect -85 -63 -81 -59
rect -101 -71 -97 -67
rect -88 -87 -84 -83
rect -52 -95 -48 -91
rect 60 -91 64 -87
rect 68 -75 72 -71
rect 76 -91 80 -87
rect 84 -75 88 -71
rect 92 -91 96 -87
rect 100 -75 104 -71
rect 129 -86 133 -82
rect -88 -103 -84 -99
rect 153 -87 157 -83
rect 161 -87 165 -83
rect 169 -87 173 -83
rect 137 -102 141 -98
rect -125 -114 -121 -110
rect -49 -130 -45 -126
rect -41 -156 -37 -152
rect -33 -156 -29 -152
rect -25 -156 -21 -152
rect 76 -147 80 -143
rect 137 -149 141 -145
rect 92 -163 96 -159
rect 145 -165 149 -161
rect 153 -149 157 -145
rect 161 -149 165 -145
rect 169 -165 173 -161
rect 177 -149 181 -145
rect 193 -165 197 -161
rect 201 -149 205 -145
rect 209 -165 213 -161
rect 231 -152 235 -148
rect -85 -172 -81 -168
rect -101 -180 -97 -176
rect 255 -153 259 -149
rect 263 -153 267 -149
rect 271 -153 275 -149
rect 239 -168 243 -164
rect 44 -184 48 -180
rect -88 -196 -84 -192
rect -52 -204 -48 -200
rect 60 -200 64 -196
rect 68 -184 72 -180
rect 76 -200 80 -196
rect 84 -184 88 -180
rect 92 -200 96 -196
rect 100 -184 104 -180
rect -88 -212 -84 -208
rect -125 -223 -121 -219
rect -49 -239 -45 -235
rect -41 -265 -37 -261
rect -33 -265 -29 -261
rect -25 -265 -21 -261
rect 76 -256 80 -252
rect 137 -258 141 -254
rect 92 -272 96 -268
rect 145 -274 149 -270
rect 153 -258 157 -254
rect 161 -258 165 -254
rect 169 -274 173 -270
rect 177 -258 181 -254
rect 193 -274 197 -270
rect 201 -258 205 -254
rect 209 -274 213 -270
rect 231 -261 235 -257
rect -85 -281 -81 -277
rect -101 -289 -97 -285
rect 255 -262 259 -258
rect 263 -262 267 -258
rect 271 -262 275 -258
rect 239 -277 243 -273
rect 44 -293 48 -289
rect -88 -305 -84 -301
rect -52 -313 -48 -309
rect 60 -309 64 -305
rect 68 -293 72 -289
rect 76 -309 80 -305
rect 84 -293 88 -289
rect 92 -309 96 -305
rect 100 -293 104 -289
rect -88 -321 -84 -317
rect -125 -332 -121 -328
rect -49 -348 -45 -344
rect -41 -374 -37 -370
rect -33 -374 -29 -370
rect -25 -374 -21 -370
rect -85 -390 -81 -386
rect -101 -398 -97 -394
rect 44 -402 48 -398
rect -88 -414 -84 -410
rect -52 -422 -48 -418
rect 60 -418 64 -414
rect 68 -402 72 -398
rect 76 -418 80 -414
rect 84 -402 88 -398
rect 92 -418 96 -414
rect 100 -402 104 -398
rect -88 -430 -84 -426
rect -125 -441 -121 -437
rect -49 -457 -45 -453
<< polysilicon >>
rect 106 -10 108 -7
rect 122 -10 124 -9
rect 82 -13 84 -10
rect 106 -22 108 -18
rect 122 -21 124 -18
rect 107 -27 108 -22
rect 106 -30 108 -27
rect 122 -30 124 -27
rect -120 -37 -118 -34
rect -36 -39 -34 -36
rect -20 -39 -18 -38
rect 82 -45 84 -33
rect 106 -37 108 -34
rect 122 -38 124 -34
rect -36 -51 -34 -47
rect -20 -50 -18 -47
rect 49 -51 51 -48
rect 57 -51 59 -47
rect -35 -56 -34 -51
rect -120 -69 -118 -57
rect -36 -59 -34 -56
rect -20 -59 -18 -56
rect -104 -66 -101 -64
rect -81 -66 -69 -64
rect -59 -66 -56 -64
rect -36 -66 -34 -63
rect -20 -67 -18 -63
rect -120 -82 -118 -79
rect -91 -90 -88 -88
rect -48 -90 -40 -88
rect -35 -90 -30 -88
rect 10 -90 13 -88
rect 82 -58 84 -55
rect 73 -71 75 -68
rect 89 -71 91 -68
rect 97 -71 99 -68
rect 158 -79 160 -76
rect 174 -79 176 -78
rect 134 -82 136 -79
rect -91 -98 -88 -96
rect -48 -98 -30 -96
rect 10 -98 13 -96
rect 49 -103 51 -91
rect 57 -103 59 -91
rect 73 -103 75 -91
rect 89 -103 91 -91
rect 97 -103 99 -91
rect 158 -91 160 -87
rect 174 -90 176 -87
rect 159 -96 160 -91
rect 158 -99 160 -96
rect 174 -99 176 -96
rect -128 -117 -125 -115
rect -45 -117 -33 -115
rect 7 -117 10 -115
rect 73 -116 75 -113
rect 134 -114 136 -102
rect 158 -106 160 -103
rect 174 -107 176 -103
rect -128 -125 -125 -123
rect -45 -125 -41 -123
rect -36 -125 -33 -123
rect 7 -125 10 -123
rect 49 -126 51 -123
rect 57 -126 59 -123
rect 89 -126 91 -123
rect 97 -125 99 -123
rect 134 -127 136 -124
rect -36 -148 -34 -145
rect -20 -148 -18 -147
rect 51 -150 54 -148
rect 64 -150 67 -148
rect 142 -145 144 -142
rect 150 -145 152 -142
rect 166 -145 168 -142
rect 182 -145 184 -142
rect 190 -145 192 -142
rect 206 -145 208 -142
rect 260 -145 262 -142
rect 276 -145 278 -144
rect 72 -150 76 -148
rect 96 -150 99 -148
rect -36 -160 -34 -156
rect -20 -159 -18 -156
rect 51 -158 54 -156
rect 64 -158 76 -156
rect 96 -158 99 -156
rect -35 -165 -34 -160
rect 236 -148 238 -145
rect -36 -168 -34 -165
rect -20 -168 -18 -165
rect -104 -175 -101 -173
rect -81 -175 -69 -173
rect -59 -175 -56 -173
rect -36 -175 -34 -172
rect -20 -176 -18 -172
rect 142 -177 144 -165
rect 150 -177 152 -165
rect 166 -177 168 -165
rect 182 -177 184 -165
rect 190 -169 192 -165
rect 190 -177 192 -174
rect 206 -177 208 -165
rect 260 -157 262 -153
rect 276 -156 278 -153
rect 261 -162 262 -157
rect 260 -165 262 -162
rect 276 -165 278 -162
rect 49 -180 51 -177
rect 57 -180 59 -177
rect 73 -180 75 -177
rect 89 -180 91 -177
rect 97 -180 99 -177
rect -91 -199 -88 -197
rect -48 -199 -40 -197
rect -35 -199 -30 -197
rect 10 -199 13 -197
rect 236 -180 238 -168
rect 260 -172 262 -169
rect 276 -173 278 -169
rect 166 -190 168 -187
rect 182 -190 184 -187
rect 190 -190 192 -187
rect 206 -190 208 -187
rect 236 -193 238 -190
rect 142 -200 144 -197
rect 150 -199 152 -197
rect -91 -207 -88 -205
rect -48 -207 -30 -205
rect 10 -207 13 -205
rect 49 -212 51 -200
rect 57 -212 59 -200
rect 73 -212 75 -200
rect 89 -212 91 -200
rect 97 -212 99 -200
rect -128 -226 -125 -224
rect -45 -226 -33 -224
rect 7 -226 10 -224
rect 49 -225 51 -222
rect 57 -225 59 -222
rect 73 -225 75 -222
rect -128 -234 -125 -232
rect -45 -234 -41 -232
rect -36 -234 -33 -232
rect 7 -234 10 -232
rect 89 -235 91 -232
rect 97 -234 99 -232
rect -36 -257 -34 -254
rect -20 -257 -18 -256
rect 51 -259 54 -257
rect 64 -259 67 -257
rect 142 -254 144 -251
rect 150 -254 152 -251
rect 166 -254 168 -251
rect 182 -254 184 -251
rect 190 -254 192 -251
rect 206 -254 208 -251
rect 260 -254 262 -251
rect 276 -254 278 -253
rect 72 -259 76 -257
rect 96 -259 99 -257
rect -36 -269 -34 -265
rect -20 -268 -18 -265
rect 51 -267 54 -265
rect 64 -267 76 -265
rect 96 -267 99 -265
rect -35 -274 -34 -269
rect 236 -257 238 -254
rect -36 -277 -34 -274
rect -20 -277 -18 -274
rect -104 -284 -101 -282
rect -81 -284 -69 -282
rect -59 -284 -56 -282
rect -36 -284 -34 -281
rect -20 -285 -18 -281
rect 142 -286 144 -274
rect 150 -286 152 -274
rect 166 -286 168 -274
rect 182 -286 184 -274
rect 190 -278 192 -274
rect 190 -286 192 -283
rect 206 -286 208 -274
rect 260 -266 262 -262
rect 276 -265 278 -262
rect 261 -271 262 -266
rect 260 -274 262 -271
rect 276 -274 278 -271
rect 49 -289 51 -286
rect 57 -289 59 -286
rect 73 -289 75 -286
rect 89 -289 91 -286
rect 97 -289 99 -286
rect -91 -308 -88 -306
rect -48 -308 -40 -306
rect -35 -308 -30 -306
rect 10 -308 13 -306
rect 236 -289 238 -277
rect 260 -281 262 -278
rect 276 -282 278 -278
rect 166 -299 168 -296
rect 182 -299 184 -296
rect 190 -299 192 -296
rect 206 -299 208 -296
rect 236 -302 238 -299
rect 142 -309 144 -306
rect 150 -308 152 -306
rect -91 -316 -88 -314
rect -48 -316 -30 -314
rect 10 -316 13 -314
rect 49 -321 51 -309
rect 57 -321 59 -309
rect 73 -321 75 -309
rect 89 -321 91 -309
rect 97 -321 99 -309
rect -128 -335 -125 -333
rect -45 -335 -33 -333
rect 7 -335 10 -333
rect 49 -334 51 -331
rect 57 -334 59 -331
rect 73 -334 75 -331
rect -128 -343 -125 -341
rect -45 -343 -41 -341
rect -36 -343 -33 -341
rect 7 -343 10 -341
rect 89 -344 91 -341
rect 97 -343 99 -341
rect -36 -366 -34 -363
rect -20 -366 -18 -365
rect -36 -378 -34 -374
rect -20 -377 -18 -374
rect -35 -383 -34 -378
rect -36 -386 -34 -383
rect -20 -386 -18 -383
rect -104 -393 -101 -391
rect -81 -393 -69 -391
rect -59 -393 -56 -391
rect -36 -393 -34 -390
rect -20 -394 -18 -390
rect 49 -398 51 -395
rect 57 -398 59 -389
rect 73 -398 75 -395
rect 89 -398 91 -395
rect 97 -398 99 -395
rect -91 -417 -88 -415
rect -48 -417 -40 -415
rect -35 -417 -30 -415
rect 10 -417 13 -415
rect -91 -425 -88 -423
rect -48 -425 -30 -423
rect 10 -425 13 -423
rect 49 -430 51 -418
rect 57 -430 59 -418
rect 73 -430 75 -418
rect 89 -430 91 -418
rect 97 -430 99 -418
rect -128 -444 -125 -442
rect -45 -444 -33 -442
rect 7 -444 10 -442
rect 49 -443 51 -440
rect 57 -443 59 -440
rect 73 -443 75 -440
rect -128 -452 -125 -450
rect -45 -452 -41 -450
rect -36 -452 -33 -450
rect 7 -452 10 -450
rect 89 -453 91 -450
rect 97 -452 99 -450
<< polycontact >>
rect 120 -9 124 -5
rect -22 -38 -18 -34
rect 78 -44 82 -40
rect 120 -42 124 -38
rect -124 -68 -120 -64
rect -74 -70 -70 -66
rect -22 -71 -18 -67
rect 172 -78 176 -74
rect 45 -96 49 -92
rect -44 -102 -40 -98
rect 69 -102 73 -98
rect 85 -101 89 -97
rect -44 -115 -40 -111
rect 130 -113 134 -109
rect 172 -111 176 -107
rect 95 -129 99 -125
rect -22 -147 -18 -143
rect 274 -144 278 -140
rect 71 -162 75 -158
rect -74 -179 -70 -175
rect 138 -170 142 -166
rect -22 -180 -18 -176
rect 162 -170 166 -166
rect 178 -170 182 -166
rect 202 -176 206 -172
rect 232 -179 236 -175
rect 274 -177 278 -173
rect 45 -205 49 -201
rect -44 -211 -40 -207
rect 69 -211 73 -207
rect 85 -210 89 -206
rect 148 -203 152 -199
rect -44 -224 -40 -220
rect 95 -238 99 -234
rect -22 -256 -18 -252
rect 274 -253 278 -249
rect 71 -271 75 -267
rect -74 -288 -70 -284
rect 138 -279 142 -275
rect -22 -289 -18 -285
rect 162 -279 166 -275
rect 178 -279 182 -275
rect 202 -285 206 -281
rect 232 -288 236 -284
rect 274 -286 278 -282
rect 45 -314 49 -310
rect -44 -320 -40 -316
rect 69 -320 73 -316
rect 85 -319 89 -315
rect 148 -312 152 -308
rect -44 -333 -40 -329
rect 95 -347 99 -343
rect -22 -365 -18 -361
rect -74 -397 -70 -393
rect -22 -398 -18 -394
rect 45 -423 49 -419
rect -44 -429 -40 -425
rect 69 -429 73 -425
rect 85 -428 89 -424
rect -44 -442 -40 -438
rect 95 -456 99 -452
<< metal1 >>
rect 96 -9 120 -6
rect 62 -17 77 -14
rect 96 -14 99 -9
rect 17 -22 41 -20
rect -131 -23 54 -22
rect -131 -25 20 -23
rect 38 -25 54 -23
rect -131 -64 -128 -25
rect -125 -31 27 -28
rect 62 -28 65 -17
rect 96 -18 101 -14
rect 96 -20 99 -18
rect 32 -31 65 -28
rect 72 -23 99 -20
rect -125 -37 -122 -31
rect -116 -37 -109 -34
rect -116 -53 -113 -37
rect -131 -67 -124 -64
rect -116 -69 -113 -57
rect -100 -67 -97 -31
rect -46 -38 -22 -35
rect 72 -36 75 -23
rect 110 -25 113 -18
rect 117 -23 120 -18
rect 117 -25 156 -23
rect 110 -26 156 -25
rect 110 -28 120 -26
rect 110 -30 113 -28
rect -46 -43 -43 -38
rect 22 -39 75 -36
rect -125 -82 -122 -79
rect -125 -85 -116 -82
rect -100 -91 -97 -71
rect -91 -46 -41 -43
rect -91 -77 -88 -46
rect -32 -54 -29 -47
rect -25 -52 -22 -47
rect 22 -52 25 -39
rect 72 -40 75 -39
rect 86 -38 89 -33
rect 117 -30 120 -28
rect 101 -38 104 -34
rect 72 -43 78 -40
rect 86 -41 120 -38
rect 86 -45 89 -41
rect -25 -54 25 -52
rect -32 -55 25 -54
rect 40 -54 44 -51
rect 48 -54 71 -51
rect -32 -57 -22 -55
rect -32 -59 -29 -57
rect -81 -62 -69 -59
rect -65 -62 -41 -59
rect -25 -59 -22 -57
rect -41 -67 -38 -63
rect 68 -65 71 -54
rect 77 -58 80 -55
rect 77 -61 112 -58
rect -74 -77 -71 -70
rect -41 -70 -22 -67
rect 68 -68 123 -65
rect 68 -71 71 -68
rect 84 -71 87 -68
rect 101 -71 104 -68
rect -62 -74 -59 -71
rect -62 -77 14 -74
rect 120 -73 123 -68
rect 120 -76 132 -73
rect -91 -80 -68 -77
rect -88 -91 -85 -87
rect -100 -94 -85 -91
rect -100 -103 -97 -94
rect -88 -99 -85 -94
rect -132 -106 -97 -103
rect -132 -110 -129 -106
rect -71 -107 -68 -80
rect -46 -83 -27 -80
rect -46 -91 -43 -83
rect -26 -86 -16 -83
rect -48 -94 -43 -91
rect -44 -107 -41 -102
rect -71 -110 -41 -107
rect -132 -113 -125 -110
rect -132 -212 -129 -113
rect -44 -111 -41 -110
rect -33 -126 -30 -114
rect -19 -126 -16 -86
rect 11 -99 14 -77
rect 129 -82 132 -76
rect 148 -78 172 -75
rect 148 -83 151 -78
rect 148 -87 153 -83
rect 148 -89 151 -87
rect 124 -90 151 -89
rect 25 -95 45 -92
rect 10 -103 14 -99
rect 61 -98 64 -91
rect 77 -98 80 -91
rect 93 -93 96 -91
rect 117 -92 151 -90
rect 117 -93 127 -92
rect 93 -96 120 -93
rect 61 -101 69 -98
rect 61 -103 64 -101
rect 77 -101 85 -98
rect 77 -103 80 -101
rect 101 -103 104 -96
rect 11 -118 14 -103
rect 48 -106 60 -103
rect 61 -112 64 -107
rect 124 -109 127 -93
rect 162 -94 165 -87
rect 169 -92 172 -87
rect 169 -94 198 -92
rect 162 -95 198 -94
rect 162 -97 172 -95
rect 162 -99 165 -97
rect 138 -107 141 -102
rect 169 -99 172 -97
rect 153 -107 156 -103
rect 124 -112 130 -109
rect 138 -110 172 -107
rect 7 -122 10 -119
rect 68 -119 71 -113
rect 138 -114 141 -110
rect 84 -119 112 -116
rect 15 -122 52 -119
rect 56 -122 84 -119
rect 117 -119 128 -116
rect 125 -120 128 -119
rect 125 -123 129 -120
rect -48 -132 -45 -130
rect -19 -129 95 -126
rect -33 -132 -29 -130
rect -48 -135 20 -132
rect 43 -137 46 -129
rect 50 -136 120 -133
rect -46 -147 -22 -144
rect 50 -145 53 -136
rect 61 -142 120 -139
rect 61 -143 64 -142
rect -46 -152 -43 -147
rect 4 -148 53 -145
rect 76 -143 80 -142
rect -91 -155 -41 -152
rect -100 -200 -97 -180
rect -91 -186 -88 -155
rect -32 -163 -29 -156
rect -25 -161 -22 -156
rect 4 -161 7 -148
rect 15 -154 54 -151
rect -25 -163 7 -161
rect -32 -164 7 -163
rect -32 -166 -22 -164
rect -32 -168 -29 -166
rect -81 -171 -69 -168
rect -65 -171 -41 -168
rect -25 -168 -22 -166
rect -41 -176 -38 -172
rect -74 -186 -71 -179
rect -41 -179 -22 -176
rect -62 -183 -59 -180
rect 11 -183 14 -156
rect 61 -159 64 -147
rect 72 -166 75 -162
rect 96 -163 103 -160
rect -62 -186 14 -183
rect -91 -189 -68 -186
rect -88 -200 -85 -196
rect -100 -203 -85 -200
rect -100 -212 -97 -203
rect -88 -208 -85 -203
rect -132 -215 -97 -212
rect -132 -219 -129 -215
rect -71 -216 -68 -189
rect -46 -192 -27 -189
rect -46 -200 -43 -192
rect -26 -195 -16 -192
rect -48 -203 -43 -200
rect -44 -216 -41 -211
rect -71 -219 -41 -216
rect -132 -222 -125 -219
rect -132 -321 -129 -222
rect -44 -220 -41 -219
rect -33 -235 -30 -223
rect -19 -235 -16 -195
rect 11 -208 14 -186
rect 21 -169 75 -166
rect 21 -200 24 -169
rect 100 -180 103 -163
rect 37 -183 44 -180
rect 48 -183 68 -180
rect 72 -183 84 -180
rect 88 -183 100 -180
rect 64 -200 68 -197
rect 25 -204 45 -201
rect 10 -212 14 -208
rect 65 -207 68 -200
rect 77 -207 80 -200
rect 93 -202 96 -200
rect 117 -200 120 -142
rect 134 -142 234 -139
rect 137 -145 140 -142
rect 154 -145 157 -142
rect 161 -145 164 -142
rect 177 -145 180 -142
rect 201 -145 204 -142
rect 231 -148 234 -142
rect 250 -144 274 -141
rect 250 -149 253 -144
rect 250 -153 255 -149
rect 250 -155 253 -153
rect 226 -158 253 -155
rect 197 -165 201 -162
rect 124 -170 138 -167
rect 146 -167 149 -165
rect 146 -170 162 -167
rect 170 -167 173 -165
rect 170 -170 178 -167
rect 154 -177 157 -170
rect 170 -177 173 -170
rect 198 -172 201 -165
rect 210 -172 213 -165
rect 226 -172 229 -158
rect 264 -160 267 -153
rect 271 -158 274 -153
rect 271 -160 292 -158
rect 264 -161 292 -160
rect 264 -163 274 -161
rect 264 -165 267 -163
rect 198 -176 202 -172
rect 210 -175 229 -172
rect 240 -173 243 -168
rect 271 -165 274 -163
rect 255 -173 258 -169
rect 198 -177 201 -176
rect 210 -177 213 -175
rect 181 -180 193 -177
rect 197 -180 201 -177
rect 226 -178 232 -175
rect 240 -176 274 -173
rect 240 -180 243 -176
rect 161 -190 164 -187
rect 186 -190 189 -187
rect 201 -190 204 -187
rect 137 -193 235 -190
rect 93 -205 109 -202
rect 65 -211 69 -207
rect 77 -210 85 -207
rect 65 -212 68 -211
rect 77 -212 80 -210
rect 101 -212 104 -205
rect 117 -203 148 -200
rect 11 -225 14 -212
rect 48 -215 60 -212
rect 64 -215 68 -212
rect 53 -225 56 -222
rect 68 -225 71 -222
rect 157 -225 160 -193
rect 11 -227 160 -225
rect 7 -231 10 -228
rect 15 -228 160 -227
rect -48 -241 -45 -239
rect -19 -238 95 -235
rect -33 -241 -29 -239
rect -48 -244 20 -241
rect 43 -246 46 -238
rect 50 -245 120 -242
rect -46 -256 -22 -253
rect 50 -254 53 -245
rect 61 -251 120 -248
rect 61 -252 64 -251
rect -46 -261 -43 -256
rect 4 -257 53 -254
rect 76 -252 80 -251
rect -91 -264 -41 -261
rect -100 -309 -97 -289
rect -91 -295 -88 -264
rect -32 -272 -29 -265
rect -25 -270 -22 -265
rect 4 -270 7 -257
rect 15 -263 54 -260
rect -25 -272 7 -270
rect -32 -273 7 -272
rect -32 -275 -22 -273
rect -32 -277 -29 -275
rect -81 -280 -69 -277
rect -65 -280 -41 -277
rect -25 -277 -22 -275
rect -41 -285 -38 -281
rect -74 -295 -71 -288
rect -41 -288 -22 -285
rect -62 -292 -59 -289
rect 11 -292 14 -265
rect 61 -268 64 -256
rect 72 -275 75 -271
rect 96 -272 103 -269
rect -62 -295 14 -292
rect -91 -298 -68 -295
rect -88 -309 -85 -305
rect -100 -312 -85 -309
rect -100 -321 -97 -312
rect -88 -317 -85 -312
rect -132 -324 -97 -321
rect -132 -328 -129 -324
rect -71 -325 -68 -298
rect -46 -301 -27 -298
rect -46 -309 -43 -301
rect -26 -304 -16 -301
rect -48 -312 -43 -309
rect -44 -325 -41 -320
rect -71 -328 -41 -325
rect -132 -331 -125 -328
rect -132 -430 -129 -331
rect -44 -329 -41 -328
rect -33 -344 -30 -332
rect -19 -344 -16 -304
rect 11 -317 14 -295
rect 21 -278 75 -275
rect 21 -309 24 -278
rect 100 -289 103 -272
rect 37 -292 44 -289
rect 48 -292 68 -289
rect 72 -292 84 -289
rect 88 -292 100 -289
rect 64 -309 68 -306
rect 25 -313 45 -310
rect 10 -321 14 -317
rect 65 -316 68 -309
rect 77 -316 80 -309
rect 93 -311 96 -309
rect 117 -309 120 -251
rect 134 -251 234 -248
rect 137 -254 140 -251
rect 154 -254 157 -251
rect 161 -254 164 -251
rect 177 -254 180 -251
rect 201 -254 204 -251
rect 231 -257 234 -251
rect 250 -253 274 -250
rect 250 -258 253 -253
rect 250 -262 255 -258
rect 250 -264 253 -262
rect 226 -267 253 -264
rect 197 -274 201 -271
rect 124 -279 138 -276
rect 146 -276 149 -274
rect 146 -279 162 -276
rect 170 -276 173 -274
rect 170 -279 178 -276
rect 154 -286 157 -279
rect 170 -286 173 -279
rect 198 -281 201 -274
rect 210 -281 213 -274
rect 226 -281 229 -267
rect 264 -269 267 -262
rect 271 -267 274 -262
rect 271 -269 288 -267
rect 264 -270 288 -269
rect 264 -272 274 -270
rect 264 -274 267 -272
rect 198 -285 202 -281
rect 210 -284 229 -281
rect 240 -282 243 -277
rect 271 -274 274 -272
rect 255 -282 258 -278
rect 198 -286 201 -285
rect 210 -286 213 -284
rect 181 -289 193 -286
rect 197 -289 201 -286
rect 226 -287 232 -284
rect 240 -285 274 -282
rect 240 -289 243 -285
rect 161 -299 164 -296
rect 186 -299 189 -296
rect 201 -299 204 -296
rect 137 -302 235 -299
rect 93 -314 109 -311
rect 65 -320 69 -316
rect 77 -319 85 -316
rect 65 -321 68 -320
rect 77 -321 80 -319
rect 101 -321 104 -314
rect 117 -312 148 -309
rect 11 -334 14 -321
rect 48 -324 60 -321
rect 64 -324 68 -321
rect 53 -334 56 -331
rect 68 -334 71 -331
rect 157 -334 160 -302
rect 11 -336 160 -334
rect 7 -340 10 -337
rect 15 -337 160 -336
rect -48 -350 -45 -348
rect -19 -347 42 -344
rect 47 -347 95 -344
rect -33 -350 -29 -348
rect -48 -353 20 -350
rect 25 -354 70 -351
rect -46 -365 -22 -362
rect -46 -370 -43 -365
rect -91 -373 -41 -370
rect -100 -418 -97 -398
rect -91 -404 -88 -373
rect -32 -381 -29 -374
rect -25 -379 -22 -374
rect 48 -379 67 -378
rect -25 -381 83 -379
rect -32 -382 51 -381
rect 64 -382 83 -381
rect -32 -384 -22 -382
rect -32 -386 -29 -384
rect -81 -389 -69 -386
rect -65 -389 -41 -386
rect -25 -386 -22 -384
rect -41 -394 -38 -390
rect -74 -404 -71 -397
rect -41 -397 -22 -394
rect 37 -395 110 -392
rect 44 -398 47 -395
rect 68 -398 71 -395
rect 84 -398 87 -395
rect 101 -398 104 -395
rect -62 -401 -59 -398
rect 11 -401 14 -398
rect -62 -404 14 -401
rect -91 -407 -68 -404
rect -88 -418 -85 -414
rect -100 -421 -85 -418
rect -100 -430 -97 -421
rect -88 -426 -85 -421
rect -132 -433 -97 -430
rect -132 -437 -129 -433
rect -71 -434 -68 -407
rect -46 -410 -27 -407
rect -46 -418 -43 -410
rect -26 -413 -16 -410
rect -48 -421 -43 -418
rect -44 -434 -41 -429
rect -71 -437 -41 -434
rect -132 -440 -125 -437
rect -132 -463 -129 -440
rect -44 -438 -41 -437
rect -33 -453 -30 -441
rect -19 -453 -16 -413
rect 11 -426 14 -404
rect 64 -418 68 -415
rect 25 -422 45 -419
rect 10 -430 14 -426
rect 65 -425 68 -418
rect 77 -425 80 -418
rect 93 -420 96 -418
rect 93 -423 115 -420
rect 65 -429 69 -425
rect 77 -428 85 -425
rect 65 -430 68 -429
rect 77 -430 80 -428
rect 11 -443 14 -430
rect 48 -433 60 -430
rect 64 -433 68 -430
rect 104 -433 107 -423
rect 53 -443 56 -440
rect 68 -443 71 -440
rect 11 -445 87 -443
rect 7 -449 10 -446
rect 15 -446 87 -445
rect -48 -459 -45 -457
rect -19 -456 95 -453
rect -33 -459 -29 -457
rect -48 -462 20 -459
<< m2contact >>
rect 54 -25 59 -20
rect -109 -39 -104 -34
rect -116 -86 -111 -81
rect 112 -62 117 -57
rect 20 -96 25 -91
rect 10 -123 15 -118
rect 112 -120 117 -115
rect 20 -137 25 -132
rect 120 -136 125 -131
rect 42 -142 47 -137
rect 10 -156 15 -151
rect 20 -205 25 -200
rect 123 -167 128 -162
rect 109 -206 114 -201
rect 10 -232 15 -227
rect 20 -246 25 -241
rect 120 -245 125 -240
rect 42 -251 47 -246
rect 10 -265 15 -260
rect 20 -314 25 -309
rect 123 -276 128 -271
rect 109 -315 114 -310
rect 10 -341 15 -336
rect 42 -347 47 -342
rect 20 -355 25 -350
rect 10 -398 15 -393
rect 20 -423 25 -418
rect 10 -450 15 -445
rect 20 -464 25 -459
<< pm12contact >>
rect 102 -27 107 -22
rect -40 -56 -35 -51
rect 56 -47 61 -42
rect -40 -92 -35 -87
rect -41 -128 -36 -123
rect 154 -96 159 -91
rect -40 -165 -35 -160
rect 67 -150 72 -145
rect -40 -201 -35 -196
rect -41 -237 -36 -232
rect 56 -177 61 -172
rect 190 -174 195 -169
rect 256 -162 261 -157
rect -40 -274 -35 -269
rect 67 -259 72 -254
rect -40 -310 -35 -305
rect -41 -346 -36 -341
rect 56 -286 61 -281
rect 190 -283 195 -278
rect 256 -271 261 -266
rect -40 -383 -35 -378
rect 56 -389 61 -384
rect -40 -419 -35 -414
rect -41 -455 -36 -450
<< pdm12contact >>
rect 125 -18 130 -13
rect -17 -47 -12 -42
rect 177 -87 182 -82
rect -17 -156 -12 -151
rect 279 -153 284 -148
rect -17 -265 -12 -260
rect 279 -262 284 -257
rect -17 -374 -12 -369
<< ndm12contact >>
rect 125 -35 130 -30
rect -17 -64 -12 -59
rect 177 -104 182 -99
rect -17 -173 -12 -168
rect 279 -170 284 -165
rect -17 -282 -12 -277
rect 279 -279 284 -274
rect -17 -391 -12 -386
<< metal2 >>
rect 126 -22 129 -18
rect 59 -23 69 -22
rect 59 -24 76 -23
rect 59 -25 102 -24
rect 66 -27 102 -25
rect 107 -25 129 -22
rect -104 -38 60 -35
rect 57 -42 60 -38
rect -16 -51 -13 -47
rect -35 -54 -13 -51
rect -116 -137 -113 -86
rect -39 -87 -36 -56
rect -16 -59 -13 -54
rect -39 -123 -36 -92
rect 11 -137 14 -123
rect 21 -132 24 -96
rect 66 -123 69 -27
rect 126 -30 129 -25
rect 113 -115 116 -62
rect 178 -91 181 -87
rect 120 -96 154 -93
rect 159 -94 181 -91
rect 66 -126 108 -123
rect 34 -132 71 -130
rect 25 -133 71 -132
rect 25 -135 37 -133
rect -116 -140 14 -137
rect 11 -151 14 -140
rect -16 -160 -13 -156
rect -35 -163 -13 -160
rect -39 -196 -36 -165
rect -16 -168 -13 -163
rect 43 -172 46 -142
rect 68 -145 71 -133
rect 105 -162 108 -126
rect 121 -131 124 -96
rect 178 -99 181 -94
rect 280 -157 283 -153
rect 221 -162 256 -159
rect 261 -160 283 -157
rect 105 -165 123 -162
rect 43 -175 56 -172
rect 110 -174 190 -171
rect -39 -232 -36 -201
rect 110 -201 113 -174
rect 11 -260 14 -232
rect 21 -241 24 -205
rect 221 -207 224 -162
rect 280 -165 283 -160
rect 121 -210 224 -207
rect 35 -241 71 -239
rect 121 -240 124 -210
rect 25 -242 71 -241
rect 25 -244 38 -242
rect -16 -269 -13 -265
rect -35 -272 -13 -269
rect -39 -305 -36 -274
rect -16 -277 -13 -272
rect 43 -281 46 -251
rect 68 -254 71 -242
rect 280 -266 283 -262
rect 221 -271 256 -268
rect 261 -269 283 -266
rect 43 -284 56 -281
rect 110 -283 190 -280
rect -39 -341 -36 -310
rect 110 -310 113 -283
rect 221 -306 224 -271
rect 280 -274 283 -269
rect -16 -378 -13 -374
rect -35 -381 -13 -378
rect -39 -414 -36 -383
rect -16 -386 -13 -381
rect 11 -393 14 -341
rect 21 -350 24 -314
rect 43 -384 46 -347
rect 43 -387 56 -384
rect -39 -450 -36 -419
rect 11 -463 14 -450
rect 21 -459 24 -423
<< m3contact >>
rect 32 -293 37 -288
<< m123contact >>
rect 27 -31 32 -26
rect 35 -55 40 -50
rect 129 -143 134 -138
rect 32 -185 37 -180
rect 129 -252 134 -247
rect 32 -396 37 -391
<< metal3 >>
rect 28 -51 31 -31
rect 28 -54 35 -51
rect 28 -139 31 -54
rect 28 -142 129 -139
rect 28 -180 31 -142
rect 28 -185 32 -180
rect 28 -248 31 -185
rect 28 -251 129 -248
rect 28 -288 31 -251
rect 28 -293 32 -288
rect 28 -391 31 -293
rect 28 -396 32 -391
use XOR  XOR_0
timestamp 1731446490
transform 1 0 567 0 1 132
box -351 -83 -274 -26
use last  last_0
timestamp 1731492129
transform 1 0 215 0 1 159
box -159 -109 -58 -45
<< labels >>
rlabel metal1 17 -243 17 -243 1 Pt1
rlabel metal1 17 -352 17 -352 1 Pt2
rlabel metal1 18 -461 18 -461 1 Pt3
rlabel metal1 18 -455 18 -455 1 G3
rlabel metal1 17 -346 17 -346 1 G2
rlabel metal1 17 -237 17 -237 1 G1
rlabel metal1 16 -381 16 -381 1 pgxor3
rlabel metal2 -37 -436 -37 -436 1 B_3
rlabel metal1 -43 -436 -43 -436 1 A_3
rlabel metal2 -38 -327 -38 -327 1 B_2
rlabel metal1 -42 -327 -42 -327 1 A_2
rlabel metal2 -38 -217 -38 -217 1 B_1
rlabel metal1 -42 -217 -42 -217 1 A_1
rlabel metal1 13 -441 13 -441 7 gnd
rlabel metal1 -131 -443 -131 -443 3 VDD
rlabel metal1 13 -332 13 -332 7 gnd
rlabel metal1 -131 -334 -131 -334 3 VDD
rlabel metal1 16 -54 16 -54 1 pgxor0
rlabel metal1 13 -114 13 -114 7 gnd
rlabel metal1 -131 -116 -131 -116 3 VDD
rlabel metal1 13 -223 13 -223 7 gnd
rlabel metal1 -131 -225 -131 -225 3 VDD
rlabel metal1 -43 -109 -43 -109 1 A_0
rlabel metal2 -38 -109 -38 -109 1 B_0
rlabel metal1 17 -134 17 -134 1 Pt0
rlabel metal1 17 -128 17 -128 1 G0
rlabel metal1 39 -203 39 -203 1 Pt1
rlabel metal1 61 -227 61 -227 1 gnd
rlabel metal1 61 -336 61 -336 1 gnd
rlabel m2contact 112 -313 112 -313 7 GPG2
rlabel metal1 39 -312 39 -312 1 Pt2
rlabel metal1 61 -445 61 -445 1 gnd
rlabel metal1 47 -394 47 -394 1 VDD
rlabel metal1 39 -421 39 -421 1 Pt3
rlabel metal1 56 -346 56 -346 1 G2
rlabel metal2 51 -386 51 -386 1 G2
rlabel metal1 111 -422 111 -422 7 GPG3
rlabel metal1 -120 -84 -120 -84 1 gnd
rlabel metal1 -123 -29 -123 -29 5 VDD
rlabel metal1 -115 -67 -115 -67 1 C0bar
rlabel metal1 -129 -66 -129 -66 3 C0
rlabel metal2 48 -37 48 -37 1 C0bar
rlabel metal1 118 -95 118 -95 1 C1
rlabel metal1 82 -60 82 -60 1 gnd
rlabel metal1 139 -25 139 -25 1 S0
rlabel metal2 52 -174 52 -174 1 G0
rlabel metal1 115 -135 115 -135 1 pgxor1
rlabel metal1 131 -74 131 -74 5 VDD
rlabel metal1 109 -118 109 -118 1 gnd
rlabel metal1 193 -94 193 -94 7 S1
rlabel metal1 101 -162 101 -162 1 VDD
rlabel metal1 6 -163 6 -163 1 pgxor1
rlabel metal1 64 -141 64 -141 1 P10
rlabel metal1 107 -204 107 -204 1 GPG1
rlabel metal2 126 -173 126 -173 1 GPG1
rlabel metal1 181 -192 181 -192 1 gnd
rlabel metal1 143 -140 143 -140 5 VDD
rlabel metal1 233 -140 233 -140 5 VDD
rlabel metal1 228 -191 228 -191 1 gnd
rlabel metal2 51 -283 51 -283 1 G1
rlabel metal1 4 -272 4 -272 1 pgxor2
rlabel metal1 101 -271 101 -271 1 VDD
rlabel metal1 181 -301 181 -301 1 gnd
rlabel metal1 143 -249 143 -249 5 VDD
rlabel metal1 233 -249 233 -249 5 VDD
rlabel metal1 228 -300 228 -300 1 gnd
rlabel metal1 126 -169 126 -169 1 C0
rlabel metal1 125 -202 125 -202 1 P10
rlabel metal1 126 -311 126 -311 1 P21
rlabel metal1 125 -278 125 -278 1 C1
rlabel metal2 125 -282 125 -282 1 GPG2
rlabel metal1 114 -244 114 -244 1 pgxor2
rlabel metal2 223 -184 223 -184 1 pgxor2
rlabel metal1 216 -173 216 -173 1 C2
rlabel metal1 290 -160 290 -160 7 S2
rlabel metal2 222 -294 222 -294 1 pgxor3
rlabel metal1 286 -269 286 -269 1 S3
<< end >>
