magic
tech scmos
timestamp 1731446490
<< nwell >>
rect -319 -29 -274 -26
rect -339 -46 -274 -29
rect -339 -61 -315 -46
<< ntransistor >>
rect -304 -56 -302 -52
rect -288 -56 -286 -52
rect -328 -77 -326 -67
<< ptransistor >>
rect -328 -55 -326 -35
rect -304 -40 -302 -32
rect -288 -40 -286 -32
<< ndiffusion >>
rect -305 -56 -304 -52
rect -302 -56 -301 -52
rect -289 -56 -288 -52
rect -286 -56 -285 -52
rect -333 -73 -328 -67
rect -329 -77 -328 -73
rect -326 -71 -325 -67
rect -326 -77 -321 -71
<< pdiffusion >>
rect -329 -39 -328 -35
rect -333 -55 -328 -39
rect -326 -51 -321 -35
rect -309 -36 -304 -32
rect -305 -40 -304 -36
rect -302 -36 -297 -32
rect -302 -40 -301 -36
rect -293 -36 -288 -32
rect -289 -40 -288 -36
rect -286 -35 -281 -32
rect -286 -40 -285 -35
rect -326 -55 -325 -51
<< ndcontact >>
rect -309 -56 -305 -52
rect -301 -56 -297 -52
rect -293 -56 -289 -52
rect -333 -77 -329 -73
rect -325 -71 -321 -67
<< pdcontact >>
rect -333 -39 -329 -35
rect -309 -40 -305 -36
rect -301 -40 -297 -36
rect -293 -40 -289 -36
rect -325 -55 -321 -51
<< polysilicon >>
rect -304 -32 -302 -29
rect -288 -32 -286 -31
rect -328 -35 -326 -32
rect -304 -44 -302 -40
rect -288 -43 -286 -40
rect -303 -49 -302 -44
rect -304 -52 -302 -49
rect -288 -52 -286 -49
rect -328 -67 -326 -55
rect -304 -59 -302 -56
rect -288 -60 -286 -56
rect -328 -80 -326 -77
<< polycontact >>
rect -290 -31 -286 -27
rect -332 -66 -328 -62
rect -290 -64 -286 -60
<< metal1 >>
rect -339 -29 -319 -26
rect -333 -35 -330 -29
rect -314 -31 -290 -28
rect -314 -36 -311 -31
rect -314 -40 -309 -36
rect -314 -42 -311 -40
rect -351 -49 -347 -46
rect -338 -45 -311 -42
rect -338 -62 -335 -45
rect -300 -47 -297 -40
rect -293 -45 -290 -40
rect -293 -47 -276 -45
rect -300 -48 -276 -47
rect -300 -50 -290 -48
rect -300 -52 -297 -50
rect -324 -60 -321 -55
rect -293 -52 -290 -50
rect -309 -60 -306 -56
rect -338 -65 -332 -62
rect -324 -63 -290 -60
rect -324 -67 -321 -63
rect -333 -80 -330 -77
rect -333 -83 -321 -80
<< m2contact >>
rect -347 -49 -342 -44
<< pm12contact >>
rect -308 -49 -303 -44
<< pdm12contact >>
rect -285 -40 -280 -35
<< ndm12contact >>
rect -285 -57 -280 -52
<< metal2 >>
rect -284 -44 -281 -40
rect -342 -49 -308 -46
rect -303 -47 -281 -44
rect -284 -52 -281 -47
<< labels >>
rlabel metal1 -331 -27 -331 -27 5 VDD
rlabel metal1 -328 -82 -328 -82 1 gnd
rlabel metal1 -350 -48 -350 -48 1 B
rlabel metal1 -336 -64 -336 -64 1 A
rlabel metal1 -277 -47 -277 -47 1 out
<< end >>
