magic
tech scmos
timestamp 1731604463
<< nwell >>
rect 71 -23 95 -11
rect 71 -31 128 -23
rect -131 -51 -107 -31
rect 59 -33 128 -31
rect -131 -63 -75 -51
rect -47 -53 -6 -33
rect 58 -43 128 -33
rect 58 -45 71 -43
rect -107 -77 -75 -63
rect 38 -65 70 -45
rect -94 -92 -36 -77
rect -94 -104 -39 -92
rect 38 -97 110 -65
rect 143 -76 188 -73
rect 123 -93 188 -76
rect -131 -136 -39 -104
rect 123 -108 147 -93
rect -47 -162 -6 -142
rect -107 -186 -75 -162
rect 70 -174 102 -137
rect 137 -151 242 -139
rect 137 -171 275 -151
rect -94 -201 -36 -186
rect -94 -213 -39 -201
rect 38 -206 110 -174
rect -131 -245 -39 -213
rect -47 -271 -6 -251
rect -107 -295 -75 -271
rect 70 -283 102 -246
rect 137 -260 242 -248
rect 137 -280 275 -260
rect -94 -310 -36 -295
rect -94 -322 -39 -310
rect 38 -315 110 -283
rect -131 -354 -39 -322
rect -47 -380 -6 -360
rect -107 -404 -75 -380
rect 70 -385 102 -355
rect 137 -373 217 -357
rect 70 -392 103 -385
rect 137 -389 248 -373
rect -94 -419 -36 -404
rect 38 -412 110 -392
rect 185 -405 248 -389
rect 185 -409 217 -405
rect -94 -431 -39 -419
rect 38 -424 124 -412
rect 111 -425 124 -424
rect 111 -431 145 -425
rect -131 -463 -39 -431
rect 112 -457 145 -431
rect 217 -441 249 -417
rect 189 -473 241 -441
<< ntransistor >>
rect -36 -63 -34 -59
rect -20 -63 -18 -59
rect -69 -66 -59 -64
rect -120 -79 -118 -69
rect -30 -90 10 -88
rect 82 -59 84 -49
rect 98 -53 100 -49
rect 114 -53 116 -49
rect -30 -98 10 -96
rect -33 -117 7 -115
rect 49 -123 51 -103
rect 57 -123 59 -103
rect 73 -113 75 -103
rect 89 -123 91 -103
rect 97 -123 99 -103
rect 158 -103 160 -99
rect 174 -103 176 -99
rect -33 -125 7 -123
rect 134 -124 136 -114
rect 54 -150 64 -148
rect 54 -158 64 -156
rect -36 -172 -34 -168
rect -20 -172 -18 -168
rect -69 -175 -59 -173
rect -30 -199 10 -197
rect 148 -197 150 -177
rect 156 -197 158 -177
rect 172 -187 174 -177
rect 188 -187 190 -177
rect 196 -187 198 -177
rect 212 -187 214 -177
rect 229 -187 231 -177
rect 245 -181 247 -177
rect 261 -181 263 -177
rect -30 -207 10 -205
rect 49 -222 51 -212
rect 57 -222 59 -212
rect 73 -222 75 -212
rect -33 -226 7 -224
rect 89 -232 91 -212
rect 97 -232 99 -212
rect -33 -234 7 -232
rect 54 -259 64 -257
rect 54 -267 64 -265
rect -36 -281 -34 -277
rect -20 -281 -18 -277
rect -69 -284 -59 -282
rect -30 -308 10 -306
rect 148 -306 150 -286
rect 156 -306 158 -286
rect 172 -296 174 -286
rect 188 -296 190 -286
rect 196 -296 198 -286
rect 212 -296 214 -286
rect 229 -296 231 -286
rect 245 -290 247 -286
rect 261 -290 263 -286
rect -30 -316 10 -314
rect 49 -331 51 -321
rect 57 -331 59 -321
rect 73 -331 75 -321
rect -33 -335 7 -333
rect 89 -341 91 -321
rect 97 -341 99 -321
rect -33 -343 7 -341
rect 54 -368 64 -366
rect 54 -376 64 -374
rect -36 -390 -34 -386
rect -20 -390 -18 -386
rect -69 -393 -59 -391
rect -30 -417 10 -415
rect 148 -415 150 -395
rect 156 -415 158 -395
rect 172 -405 174 -395
rect 257 -386 277 -384
rect 257 -394 277 -392
rect -30 -425 10 -423
rect 49 -440 51 -430
rect 57 -440 59 -430
rect 73 -440 75 -430
rect -33 -444 7 -442
rect 89 -450 91 -430
rect 97 -450 99 -430
rect 196 -435 198 -415
rect 204 -435 206 -415
rect 255 -430 265 -428
rect 156 -438 176 -436
rect 156 -446 176 -444
rect -33 -452 7 -450
rect 247 -454 267 -452
rect 247 -462 267 -460
<< ptransistor >>
rect -120 -57 -118 -37
rect 82 -37 84 -17
rect 98 -37 100 -29
rect 114 -37 116 -29
rect -36 -47 -34 -39
rect -20 -47 -18 -39
rect -101 -66 -81 -64
rect -88 -90 -48 -88
rect 49 -91 51 -51
rect 57 -91 59 -51
rect 73 -91 75 -71
rect 89 -91 91 -71
rect 97 -91 99 -71
rect -88 -98 -48 -96
rect 134 -102 136 -82
rect 158 -87 160 -79
rect 174 -87 176 -79
rect -125 -117 -45 -115
rect -125 -125 -45 -123
rect -36 -156 -34 -148
rect -20 -156 -18 -148
rect 76 -150 96 -148
rect 76 -158 96 -156
rect 148 -165 150 -145
rect 156 -165 158 -145
rect 172 -165 174 -145
rect 188 -165 190 -145
rect 196 -165 198 -145
rect 212 -165 214 -145
rect 229 -165 231 -145
rect 245 -165 247 -157
rect 261 -165 263 -157
rect -101 -175 -81 -173
rect -88 -199 -48 -197
rect 49 -200 51 -180
rect 57 -200 59 -180
rect 73 -200 75 -180
rect 89 -200 91 -180
rect 97 -200 99 -180
rect -88 -207 -48 -205
rect -125 -226 -45 -224
rect -125 -234 -45 -232
rect -36 -265 -34 -257
rect -20 -265 -18 -257
rect 76 -259 96 -257
rect 76 -267 96 -265
rect 148 -274 150 -254
rect 156 -274 158 -254
rect 172 -274 174 -254
rect 188 -274 190 -254
rect 196 -274 198 -254
rect 212 -274 214 -254
rect 229 -274 231 -254
rect 245 -274 247 -266
rect 261 -274 263 -266
rect -101 -284 -81 -282
rect -88 -308 -48 -306
rect 49 -309 51 -289
rect 57 -309 59 -289
rect 73 -309 75 -289
rect 89 -309 91 -289
rect 97 -309 99 -289
rect -88 -316 -48 -314
rect -125 -335 -45 -333
rect -125 -343 -45 -341
rect -36 -374 -34 -366
rect -20 -374 -18 -366
rect 76 -368 96 -366
rect 76 -376 96 -374
rect 148 -383 150 -363
rect 156 -383 158 -363
rect 172 -383 174 -363
rect -101 -393 -81 -391
rect -88 -417 -48 -415
rect 49 -418 51 -398
rect 57 -418 59 -398
rect 73 -418 75 -398
rect 89 -418 91 -398
rect 97 -418 99 -398
rect 196 -403 198 -363
rect 204 -403 206 -363
rect 219 -386 239 -384
rect 219 -394 239 -392
rect -88 -425 -48 -423
rect -125 -444 -45 -442
rect 223 -430 243 -428
rect 118 -438 138 -436
rect 118 -446 138 -444
rect -125 -452 -45 -450
rect 195 -454 235 -452
rect 195 -462 235 -460
<< ndiffusion >>
rect -65 -63 -59 -59
rect -37 -63 -36 -59
rect -34 -63 -33 -59
rect -21 -63 -20 -59
rect -18 -63 -17 -59
rect -69 -64 -59 -63
rect -125 -75 -120 -69
rect -121 -79 -120 -75
rect -118 -73 -117 -69
rect -69 -67 -59 -66
rect -69 -71 -63 -67
rect -118 -79 -113 -73
rect -26 -87 10 -83
rect -30 -88 10 -87
rect -30 -96 10 -90
rect 77 -54 82 -49
rect 81 -59 82 -54
rect 84 -53 85 -49
rect 97 -53 98 -49
rect 100 -53 101 -49
rect 113 -53 114 -49
rect 116 -53 117 -49
rect 84 -59 89 -53
rect -30 -99 10 -98
rect -30 -103 6 -99
rect 48 -107 49 -103
rect -29 -114 7 -110
rect -33 -115 7 -114
rect -33 -118 7 -117
rect -33 -122 3 -118
rect -33 -123 7 -122
rect 44 -123 49 -107
rect 51 -119 57 -103
rect 51 -123 52 -119
rect 56 -123 57 -119
rect 59 -107 60 -103
rect 59 -123 64 -107
rect 68 -109 73 -103
rect 72 -113 73 -109
rect 75 -107 76 -103
rect 75 -113 80 -107
rect 84 -119 89 -103
rect 88 -123 89 -119
rect 91 -123 97 -103
rect 99 -107 100 -103
rect 99 -123 104 -107
rect 157 -103 158 -99
rect 160 -103 161 -99
rect 173 -103 174 -99
rect 176 -103 177 -99
rect 129 -120 134 -114
rect -33 -126 7 -125
rect 133 -124 134 -120
rect 136 -118 137 -114
rect 136 -124 141 -118
rect -29 -130 7 -126
rect 54 -147 60 -143
rect 54 -148 64 -147
rect 54 -151 64 -150
rect 58 -155 64 -151
rect 54 -156 64 -155
rect 54 -159 64 -158
rect 54 -163 60 -159
rect -65 -172 -59 -168
rect -37 -172 -36 -168
rect -34 -172 -33 -168
rect -21 -172 -20 -168
rect -18 -172 -17 -168
rect -69 -173 -59 -172
rect -69 -176 -59 -175
rect -69 -180 -63 -176
rect -26 -196 10 -192
rect -30 -197 10 -196
rect -30 -205 10 -199
rect 143 -193 148 -177
rect 147 -197 148 -193
rect 150 -197 156 -177
rect 158 -181 159 -177
rect 158 -197 163 -181
rect 167 -183 172 -177
rect 171 -187 172 -183
rect 174 -181 175 -177
rect 174 -187 179 -181
rect 187 -181 188 -177
rect 183 -187 188 -181
rect 190 -183 196 -177
rect 190 -187 191 -183
rect 195 -187 196 -183
rect 198 -181 199 -177
rect 198 -187 203 -181
rect 207 -183 212 -177
rect 211 -187 212 -183
rect 214 -181 215 -177
rect 214 -187 219 -181
rect 224 -183 229 -177
rect 228 -187 229 -183
rect 231 -181 232 -177
rect 244 -181 245 -177
rect 247 -181 248 -177
rect 260 -181 261 -177
rect 263 -181 264 -177
rect 231 -187 236 -181
rect -30 -208 10 -207
rect -30 -212 6 -208
rect 48 -216 49 -212
rect -29 -223 7 -219
rect 44 -222 49 -216
rect 51 -218 57 -212
rect 51 -222 52 -218
rect 56 -222 57 -218
rect 59 -216 60 -212
rect 59 -222 64 -216
rect 68 -218 73 -212
rect 72 -222 73 -218
rect 75 -216 76 -212
rect 75 -222 80 -216
rect -33 -224 7 -223
rect -33 -227 7 -226
rect -33 -231 3 -227
rect -33 -232 7 -231
rect 84 -228 89 -212
rect 88 -232 89 -228
rect 91 -232 97 -212
rect 99 -216 100 -212
rect 99 -232 104 -216
rect -33 -235 7 -234
rect -29 -239 7 -235
rect 54 -256 60 -252
rect 54 -257 64 -256
rect 54 -260 64 -259
rect 58 -264 64 -260
rect 54 -265 64 -264
rect 54 -268 64 -267
rect 54 -272 60 -268
rect -65 -281 -59 -277
rect -37 -281 -36 -277
rect -34 -281 -33 -277
rect -21 -281 -20 -277
rect -18 -281 -17 -277
rect -69 -282 -59 -281
rect -69 -285 -59 -284
rect -69 -289 -63 -285
rect -26 -305 10 -301
rect -30 -306 10 -305
rect -30 -314 10 -308
rect 143 -302 148 -286
rect 147 -306 148 -302
rect 150 -306 156 -286
rect 158 -290 159 -286
rect 158 -306 163 -290
rect 167 -292 172 -286
rect 171 -296 172 -292
rect 174 -290 175 -286
rect 174 -296 179 -290
rect 187 -290 188 -286
rect 183 -296 188 -290
rect 190 -292 196 -286
rect 190 -296 191 -292
rect 195 -296 196 -292
rect 198 -290 199 -286
rect 198 -296 203 -290
rect 207 -292 212 -286
rect 211 -296 212 -292
rect 214 -290 215 -286
rect 214 -296 219 -290
rect 224 -292 229 -286
rect 228 -296 229 -292
rect 231 -290 232 -286
rect 244 -290 245 -286
rect 247 -290 248 -286
rect 260 -290 261 -286
rect 263 -290 264 -286
rect 231 -296 236 -290
rect -30 -317 10 -316
rect -30 -321 6 -317
rect 48 -325 49 -321
rect -29 -332 7 -328
rect 44 -331 49 -325
rect 51 -327 57 -321
rect 51 -331 52 -327
rect 56 -331 57 -327
rect 59 -325 60 -321
rect 59 -331 64 -325
rect 68 -327 73 -321
rect 72 -331 73 -327
rect 75 -325 76 -321
rect 75 -331 80 -325
rect -33 -333 7 -332
rect -33 -336 7 -335
rect -33 -340 3 -336
rect -33 -341 7 -340
rect 84 -337 89 -321
rect 88 -341 89 -337
rect 91 -341 97 -321
rect 99 -325 100 -321
rect 99 -341 104 -325
rect -33 -344 7 -343
rect -29 -348 7 -344
rect 54 -365 60 -361
rect 54 -366 64 -365
rect 54 -369 64 -368
rect 58 -373 64 -369
rect 54 -374 64 -373
rect 54 -377 64 -376
rect 54 -381 60 -377
rect -65 -390 -59 -386
rect -37 -390 -36 -386
rect -34 -390 -33 -386
rect -21 -390 -20 -386
rect -18 -390 -17 -386
rect -69 -391 -59 -390
rect -69 -394 -59 -393
rect -69 -398 -63 -394
rect -26 -414 10 -410
rect -30 -415 10 -414
rect -30 -423 10 -417
rect 143 -411 148 -395
rect 147 -415 148 -411
rect 150 -415 156 -395
rect 158 -399 159 -395
rect 158 -415 163 -399
rect 167 -401 172 -395
rect 171 -405 172 -401
rect 174 -399 175 -395
rect 174 -405 179 -399
rect 261 -383 277 -379
rect 257 -384 277 -383
rect 257 -392 277 -386
rect 257 -395 277 -394
rect 257 -399 273 -395
rect -30 -426 10 -425
rect -30 -430 6 -426
rect 195 -419 196 -415
rect 48 -434 49 -430
rect -29 -441 7 -437
rect 44 -440 49 -434
rect 51 -436 57 -430
rect 51 -440 52 -436
rect 56 -440 57 -436
rect 59 -434 60 -430
rect 59 -440 64 -434
rect 68 -436 73 -430
rect 72 -440 73 -436
rect 75 -434 76 -430
rect 75 -440 80 -434
rect -33 -442 7 -441
rect -33 -445 7 -444
rect -33 -449 3 -445
rect -33 -450 7 -449
rect 84 -446 89 -430
rect 88 -450 89 -446
rect 91 -450 97 -430
rect 99 -434 100 -430
rect 99 -450 104 -434
rect 156 -435 172 -431
rect 191 -435 196 -419
rect 198 -431 204 -415
rect 198 -435 199 -431
rect 203 -435 204 -431
rect 206 -419 207 -415
rect 206 -435 211 -419
rect 259 -427 265 -423
rect 255 -428 265 -427
rect 255 -431 265 -430
rect 255 -435 261 -431
rect 156 -436 176 -435
rect 156 -444 176 -438
rect -33 -453 7 -452
rect 156 -447 176 -446
rect 160 -451 176 -447
rect -29 -457 7 -453
rect 251 -451 267 -447
rect 247 -452 267 -451
rect 247 -455 267 -454
rect 247 -459 263 -455
rect 247 -460 267 -459
rect 247 -463 267 -462
rect 251 -467 267 -463
<< pdiffusion >>
rect 81 -21 82 -17
rect -121 -41 -120 -37
rect -125 -57 -120 -41
rect -118 -53 -113 -37
rect 77 -37 82 -21
rect 84 -33 89 -17
rect 84 -37 85 -33
rect 93 -33 98 -29
rect 97 -37 98 -33
rect 100 -33 105 -29
rect 100 -37 101 -33
rect 109 -33 114 -29
rect 113 -37 114 -33
rect 116 -32 121 -29
rect 116 -37 117 -32
rect -41 -43 -36 -39
rect -37 -47 -36 -43
rect -34 -43 -29 -39
rect -34 -47 -33 -43
rect -25 -43 -20 -39
rect -21 -47 -20 -43
rect -18 -42 -13 -39
rect -18 -47 -17 -42
rect -118 -57 -117 -53
rect 48 -55 49 -51
rect -101 -63 -85 -59
rect -101 -64 -81 -63
rect -101 -67 -81 -66
rect -97 -71 -81 -67
rect -84 -87 -48 -83
rect -88 -88 -48 -87
rect -88 -91 -48 -90
rect -88 -95 -52 -91
rect -88 -96 -48 -95
rect 44 -91 49 -55
rect 51 -91 57 -51
rect 59 -87 64 -51
rect 59 -91 60 -87
rect 72 -75 73 -71
rect 68 -91 73 -75
rect 75 -87 80 -71
rect 75 -91 76 -87
rect 88 -75 89 -71
rect 84 -91 89 -75
rect 91 -87 97 -71
rect 91 -91 92 -87
rect 96 -91 97 -87
rect 99 -75 100 -71
rect 99 -91 104 -75
rect 133 -86 134 -82
rect -88 -99 -48 -98
rect -84 -103 -48 -99
rect 129 -102 134 -86
rect 136 -98 141 -82
rect 153 -83 158 -79
rect 157 -87 158 -83
rect 160 -83 165 -79
rect 160 -87 161 -83
rect 169 -83 174 -79
rect 173 -87 174 -83
rect 176 -82 181 -79
rect 176 -87 177 -82
rect 136 -102 137 -98
rect -121 -114 -45 -110
rect -125 -115 -45 -114
rect -125 -123 -45 -117
rect -125 -126 -45 -125
rect -125 -130 -49 -126
rect -41 -152 -36 -148
rect -37 -156 -36 -152
rect -34 -152 -29 -148
rect -34 -156 -33 -152
rect -25 -152 -20 -148
rect -21 -156 -20 -152
rect -18 -151 -13 -148
rect 80 -147 96 -143
rect 76 -148 96 -147
rect 147 -149 148 -145
rect -18 -156 -17 -151
rect 76 -156 96 -150
rect 76 -159 96 -158
rect 76 -163 92 -159
rect 143 -165 148 -149
rect 150 -161 156 -145
rect 150 -165 151 -161
rect 155 -165 156 -161
rect 158 -149 159 -145
rect 158 -165 163 -149
rect 171 -149 172 -145
rect 167 -165 172 -149
rect 174 -161 179 -145
rect 174 -165 175 -161
rect 187 -149 188 -145
rect 183 -165 188 -149
rect 190 -165 196 -145
rect 198 -161 203 -145
rect 198 -165 199 -161
rect 211 -149 212 -145
rect 207 -165 212 -149
rect 214 -161 219 -145
rect 214 -165 215 -161
rect 228 -149 229 -145
rect 224 -165 229 -149
rect 231 -161 236 -145
rect 231 -165 232 -161
rect 240 -161 245 -157
rect 244 -165 245 -161
rect 247 -161 252 -157
rect 247 -165 248 -161
rect 256 -161 261 -157
rect 260 -165 261 -161
rect 263 -160 268 -157
rect 263 -165 264 -160
rect -101 -172 -85 -168
rect -101 -173 -81 -172
rect -101 -176 -81 -175
rect -97 -180 -81 -176
rect 48 -184 49 -180
rect -84 -196 -48 -192
rect -88 -197 -48 -196
rect -88 -200 -48 -199
rect -88 -204 -52 -200
rect -88 -205 -48 -204
rect 44 -200 49 -184
rect 51 -200 57 -180
rect 59 -196 64 -180
rect 59 -200 60 -196
rect 72 -184 73 -180
rect 68 -200 73 -184
rect 75 -196 80 -180
rect 75 -200 76 -196
rect 88 -184 89 -180
rect 84 -200 89 -184
rect 91 -196 97 -180
rect 91 -200 92 -196
rect 96 -200 97 -196
rect 99 -184 100 -180
rect 99 -200 104 -184
rect -88 -208 -48 -207
rect -84 -212 -48 -208
rect -121 -223 -45 -219
rect -125 -224 -45 -223
rect -125 -232 -45 -226
rect -125 -235 -45 -234
rect -125 -239 -49 -235
rect -41 -261 -36 -257
rect -37 -265 -36 -261
rect -34 -261 -29 -257
rect -34 -265 -33 -261
rect -25 -261 -20 -257
rect -21 -265 -20 -261
rect -18 -260 -13 -257
rect 80 -256 96 -252
rect 76 -257 96 -256
rect 147 -258 148 -254
rect -18 -265 -17 -260
rect 76 -265 96 -259
rect 76 -268 96 -267
rect 76 -272 92 -268
rect 143 -274 148 -258
rect 150 -270 156 -254
rect 150 -274 151 -270
rect 155 -274 156 -270
rect 158 -258 159 -254
rect 158 -274 163 -258
rect 171 -258 172 -254
rect 167 -274 172 -258
rect 174 -270 179 -254
rect 174 -274 175 -270
rect 187 -258 188 -254
rect 183 -274 188 -258
rect 190 -274 196 -254
rect 198 -270 203 -254
rect 198 -274 199 -270
rect 211 -258 212 -254
rect 207 -274 212 -258
rect 214 -270 219 -254
rect 214 -274 215 -270
rect 228 -258 229 -254
rect 224 -274 229 -258
rect 231 -270 236 -254
rect 231 -274 232 -270
rect 240 -270 245 -266
rect 244 -274 245 -270
rect 247 -270 252 -266
rect 247 -274 248 -270
rect 256 -270 261 -266
rect 260 -274 261 -270
rect 263 -269 268 -266
rect 263 -274 264 -269
rect -101 -281 -85 -277
rect -101 -282 -81 -281
rect -101 -285 -81 -284
rect -97 -289 -81 -285
rect 48 -293 49 -289
rect -84 -305 -48 -301
rect -88 -306 -48 -305
rect -88 -309 -48 -308
rect -88 -313 -52 -309
rect -88 -314 -48 -313
rect 44 -309 49 -293
rect 51 -309 57 -289
rect 59 -305 64 -289
rect 59 -309 60 -305
rect 72 -293 73 -289
rect 68 -309 73 -293
rect 75 -305 80 -289
rect 75 -309 76 -305
rect 88 -293 89 -289
rect 84 -309 89 -293
rect 91 -305 97 -289
rect 91 -309 92 -305
rect 96 -309 97 -305
rect 99 -293 100 -289
rect 99 -309 104 -293
rect -88 -317 -48 -316
rect -84 -321 -48 -317
rect -121 -332 -45 -328
rect -125 -333 -45 -332
rect -125 -341 -45 -335
rect -125 -344 -45 -343
rect -125 -348 -49 -344
rect -41 -370 -36 -366
rect -37 -374 -36 -370
rect -34 -370 -29 -366
rect -34 -374 -33 -370
rect -25 -370 -20 -366
rect -21 -374 -20 -370
rect -18 -369 -13 -366
rect 80 -365 96 -361
rect 76 -366 96 -365
rect 147 -367 148 -363
rect -18 -374 -17 -369
rect 76 -374 96 -368
rect 76 -377 96 -376
rect 76 -381 92 -377
rect 143 -383 148 -367
rect 150 -379 156 -363
rect 150 -383 151 -379
rect 155 -383 156 -379
rect 158 -367 159 -363
rect 158 -383 163 -367
rect 171 -367 172 -363
rect 167 -383 172 -367
rect 174 -379 179 -363
rect 174 -383 175 -379
rect 195 -367 196 -363
rect -101 -390 -85 -386
rect -101 -391 -81 -390
rect -101 -394 -81 -393
rect -97 -398 -81 -394
rect 48 -402 49 -398
rect -84 -414 -48 -410
rect -88 -415 -48 -414
rect -88 -418 -48 -417
rect -88 -422 -52 -418
rect -88 -423 -48 -422
rect 44 -418 49 -402
rect 51 -418 57 -398
rect 59 -414 64 -398
rect 59 -418 60 -414
rect 72 -402 73 -398
rect 68 -418 73 -402
rect 75 -414 80 -398
rect 75 -418 76 -414
rect 88 -402 89 -398
rect 84 -418 89 -402
rect 91 -414 97 -398
rect 91 -418 92 -414
rect 96 -418 97 -414
rect 99 -402 100 -398
rect 99 -418 104 -402
rect 191 -403 196 -367
rect 198 -403 204 -363
rect 206 -399 211 -363
rect 223 -383 239 -379
rect 219 -384 239 -383
rect 219 -387 239 -386
rect 219 -391 235 -387
rect 219 -392 239 -391
rect 219 -395 239 -394
rect 223 -399 239 -395
rect 206 -403 207 -399
rect -88 -426 -48 -425
rect -84 -430 -48 -426
rect -121 -441 -45 -437
rect -125 -442 -45 -441
rect -125 -450 -45 -444
rect 122 -435 138 -431
rect 118 -436 138 -435
rect 223 -427 239 -423
rect 223 -428 243 -427
rect 223 -431 243 -430
rect 227 -435 243 -431
rect 118 -439 138 -438
rect 118 -443 134 -439
rect 118 -444 138 -443
rect 118 -447 138 -446
rect -125 -453 -45 -452
rect -125 -457 -49 -453
rect 122 -451 138 -447
rect 195 -451 231 -447
rect 195 -452 235 -451
rect 195 -460 235 -454
rect 195 -463 235 -462
rect 199 -467 235 -463
<< ndcontact >>
rect -69 -63 -65 -59
rect -41 -63 -37 -59
rect -33 -63 -29 -59
rect -25 -63 -21 -59
rect -125 -79 -121 -75
rect -117 -73 -113 -69
rect -63 -71 -59 -67
rect -30 -87 -26 -83
rect 85 -53 89 -49
rect 93 -53 97 -49
rect 101 -53 105 -49
rect 109 -53 113 -49
rect 6 -103 10 -99
rect 44 -107 48 -103
rect -33 -114 -29 -110
rect 3 -122 7 -118
rect 52 -123 56 -119
rect 60 -107 64 -103
rect 68 -113 72 -109
rect 76 -107 80 -103
rect 84 -123 88 -119
rect 100 -107 104 -103
rect 153 -103 157 -99
rect 161 -103 165 -99
rect 169 -103 173 -99
rect 129 -124 133 -120
rect 137 -118 141 -114
rect -33 -130 -29 -126
rect 60 -147 64 -143
rect 54 -155 58 -151
rect 60 -163 64 -159
rect -69 -172 -65 -168
rect -41 -172 -37 -168
rect -33 -172 -29 -168
rect -25 -172 -21 -168
rect -63 -180 -59 -176
rect -30 -196 -26 -192
rect 143 -197 147 -193
rect 159 -181 163 -177
rect 167 -187 171 -183
rect 175 -181 179 -177
rect 183 -181 187 -177
rect 191 -187 195 -183
rect 199 -181 203 -177
rect 207 -187 211 -183
rect 215 -181 219 -177
rect 224 -187 228 -183
rect 232 -181 236 -177
rect 240 -181 244 -177
rect 248 -181 252 -177
rect 256 -181 260 -177
rect 6 -212 10 -208
rect 44 -216 48 -212
rect -33 -223 -29 -219
rect 52 -222 56 -218
rect 60 -216 64 -212
rect 68 -222 72 -218
rect 76 -216 80 -212
rect 3 -231 7 -227
rect 84 -232 88 -228
rect 100 -216 104 -212
rect -33 -239 -29 -235
rect 60 -256 64 -252
rect 54 -264 58 -260
rect 60 -272 64 -268
rect -69 -281 -65 -277
rect -41 -281 -37 -277
rect -33 -281 -29 -277
rect -25 -281 -21 -277
rect -63 -289 -59 -285
rect -30 -305 -26 -301
rect 143 -306 147 -302
rect 159 -290 163 -286
rect 167 -296 171 -292
rect 175 -290 179 -286
rect 183 -290 187 -286
rect 191 -296 195 -292
rect 199 -290 203 -286
rect 207 -296 211 -292
rect 215 -290 219 -286
rect 224 -296 228 -292
rect 232 -290 236 -286
rect 240 -290 244 -286
rect 248 -290 252 -286
rect 256 -290 260 -286
rect 6 -321 10 -317
rect 44 -325 48 -321
rect -33 -332 -29 -328
rect 52 -331 56 -327
rect 60 -325 64 -321
rect 68 -331 72 -327
rect 76 -325 80 -321
rect 3 -340 7 -336
rect 84 -341 88 -337
rect 100 -325 104 -321
rect -33 -348 -29 -344
rect 60 -365 64 -361
rect 54 -373 58 -369
rect 60 -381 64 -377
rect -69 -390 -65 -386
rect -41 -390 -37 -386
rect -33 -390 -29 -386
rect -25 -390 -21 -386
rect -63 -398 -59 -394
rect -30 -414 -26 -410
rect 143 -415 147 -411
rect 159 -399 163 -395
rect 167 -405 171 -401
rect 175 -399 179 -395
rect 257 -383 261 -379
rect 273 -399 277 -395
rect 6 -430 10 -426
rect 191 -419 195 -415
rect 44 -434 48 -430
rect -33 -441 -29 -437
rect 52 -440 56 -436
rect 60 -434 64 -430
rect 68 -440 72 -436
rect 76 -434 80 -430
rect 3 -449 7 -445
rect 84 -450 88 -446
rect 100 -434 104 -430
rect 172 -435 176 -431
rect 199 -435 203 -431
rect 207 -419 211 -415
rect 255 -427 259 -423
rect 261 -435 265 -431
rect 156 -451 160 -447
rect -33 -457 -29 -453
rect 247 -451 251 -447
rect 263 -459 267 -455
rect 247 -467 251 -463
<< pdcontact >>
rect 77 -21 81 -17
rect -125 -41 -121 -37
rect 85 -37 89 -33
rect 93 -37 97 -33
rect 101 -37 105 -33
rect 109 -37 113 -33
rect -41 -47 -37 -43
rect -33 -47 -29 -43
rect -25 -47 -21 -43
rect -117 -57 -113 -53
rect 44 -55 48 -51
rect -85 -63 -81 -59
rect -101 -71 -97 -67
rect -88 -87 -84 -83
rect -52 -95 -48 -91
rect 60 -91 64 -87
rect 68 -75 72 -71
rect 76 -91 80 -87
rect 84 -75 88 -71
rect 92 -91 96 -87
rect 100 -75 104 -71
rect 129 -86 133 -82
rect -88 -103 -84 -99
rect 153 -87 157 -83
rect 161 -87 165 -83
rect 169 -87 173 -83
rect 137 -102 141 -98
rect -125 -114 -121 -110
rect -49 -130 -45 -126
rect -41 -156 -37 -152
rect -33 -156 -29 -152
rect -25 -156 -21 -152
rect 76 -147 80 -143
rect 143 -149 147 -145
rect 92 -163 96 -159
rect 151 -165 155 -161
rect 159 -149 163 -145
rect 167 -149 171 -145
rect 175 -165 179 -161
rect 183 -149 187 -145
rect 199 -165 203 -161
rect 207 -149 211 -145
rect 215 -165 219 -161
rect 224 -149 228 -145
rect 232 -165 236 -161
rect 240 -165 244 -161
rect 248 -165 252 -161
rect 256 -165 260 -161
rect -85 -172 -81 -168
rect -101 -180 -97 -176
rect 44 -184 48 -180
rect -88 -196 -84 -192
rect -52 -204 -48 -200
rect 60 -200 64 -196
rect 68 -184 72 -180
rect 76 -200 80 -196
rect 84 -184 88 -180
rect 92 -200 96 -196
rect 100 -184 104 -180
rect -88 -212 -84 -208
rect -125 -223 -121 -219
rect -49 -239 -45 -235
rect -41 -265 -37 -261
rect -33 -265 -29 -261
rect -25 -265 -21 -261
rect 76 -256 80 -252
rect 143 -258 147 -254
rect 92 -272 96 -268
rect 151 -274 155 -270
rect 159 -258 163 -254
rect 167 -258 171 -254
rect 175 -274 179 -270
rect 183 -258 187 -254
rect 199 -274 203 -270
rect 207 -258 211 -254
rect 215 -274 219 -270
rect 224 -258 228 -254
rect 232 -274 236 -270
rect 240 -274 244 -270
rect 248 -274 252 -270
rect 256 -274 260 -270
rect -85 -281 -81 -277
rect -101 -289 -97 -285
rect 44 -293 48 -289
rect -88 -305 -84 -301
rect -52 -313 -48 -309
rect 60 -309 64 -305
rect 68 -293 72 -289
rect 76 -309 80 -305
rect 84 -293 88 -289
rect 92 -309 96 -305
rect 100 -293 104 -289
rect -88 -321 -84 -317
rect -125 -332 -121 -328
rect -49 -348 -45 -344
rect -41 -374 -37 -370
rect -33 -374 -29 -370
rect -25 -374 -21 -370
rect 76 -365 80 -361
rect 143 -367 147 -363
rect 92 -381 96 -377
rect 151 -383 155 -379
rect 159 -367 163 -363
rect 167 -367 171 -363
rect 175 -383 179 -379
rect 191 -367 195 -363
rect -85 -390 -81 -386
rect -101 -398 -97 -394
rect 44 -402 48 -398
rect -88 -414 -84 -410
rect -52 -422 -48 -418
rect 60 -418 64 -414
rect 68 -402 72 -398
rect 76 -418 80 -414
rect 84 -402 88 -398
rect 92 -418 96 -414
rect 100 -402 104 -398
rect 219 -383 223 -379
rect 235 -391 239 -387
rect 219 -399 223 -395
rect 207 -403 211 -399
rect -88 -430 -84 -426
rect -125 -441 -121 -437
rect 118 -435 122 -431
rect 239 -427 243 -423
rect 223 -435 227 -431
rect 134 -443 138 -439
rect -49 -457 -45 -453
rect 118 -451 122 -447
rect 231 -451 235 -447
rect 195 -467 199 -463
<< polysilicon >>
rect 82 -17 84 -14
rect -120 -37 -118 -34
rect -36 -39 -34 -36
rect 98 -29 100 -26
rect 114 -29 116 -28
rect -20 -39 -18 -38
rect -36 -51 -34 -47
rect -20 -50 -18 -47
rect 49 -51 51 -48
rect 57 -51 59 -47
rect 82 -49 84 -37
rect 98 -49 100 -37
rect 114 -40 116 -37
rect 114 -49 116 -46
rect -35 -56 -34 -51
rect -120 -69 -118 -57
rect -36 -59 -34 -56
rect -20 -59 -18 -56
rect -104 -66 -101 -64
rect -81 -66 -69 -64
rect -59 -66 -56 -64
rect -36 -66 -34 -63
rect -20 -67 -18 -63
rect -120 -82 -118 -79
rect -91 -90 -88 -88
rect -48 -90 -40 -88
rect -35 -90 -30 -88
rect 10 -90 13 -88
rect 98 -56 100 -53
rect 114 -57 116 -53
rect 82 -62 84 -59
rect 73 -71 75 -68
rect 89 -71 91 -68
rect 97 -71 99 -68
rect 158 -79 160 -76
rect 174 -79 176 -78
rect 134 -82 136 -79
rect -91 -98 -88 -96
rect -48 -98 -30 -96
rect 10 -98 13 -96
rect 49 -103 51 -91
rect 57 -103 59 -91
rect 73 -103 75 -91
rect 89 -103 91 -91
rect 97 -103 99 -91
rect 158 -91 160 -87
rect 174 -90 176 -87
rect 159 -96 160 -91
rect 158 -99 160 -96
rect 174 -99 176 -96
rect -128 -117 -125 -115
rect -45 -117 -33 -115
rect 7 -117 10 -115
rect 73 -116 75 -113
rect 134 -114 136 -102
rect 158 -106 160 -103
rect 174 -107 176 -103
rect -128 -125 -125 -123
rect -45 -125 -41 -123
rect -36 -125 -33 -123
rect 7 -125 10 -123
rect 49 -126 51 -123
rect 57 -126 59 -123
rect 89 -126 91 -123
rect 97 -125 99 -123
rect 134 -127 136 -124
rect -36 -148 -34 -145
rect -20 -148 -18 -147
rect 51 -150 54 -148
rect 64 -150 67 -148
rect 148 -145 150 -142
rect 156 -145 158 -142
rect 172 -145 174 -142
rect 188 -145 190 -142
rect 196 -145 198 -142
rect 212 -145 214 -142
rect 229 -145 231 -142
rect 72 -150 76 -148
rect 96 -150 99 -148
rect -36 -160 -34 -156
rect -20 -159 -18 -156
rect 51 -158 54 -156
rect 64 -158 76 -156
rect 96 -158 99 -156
rect -35 -165 -34 -160
rect 245 -157 247 -154
rect 261 -157 263 -156
rect -36 -168 -34 -165
rect -20 -168 -18 -165
rect -104 -175 -101 -173
rect -81 -175 -69 -173
rect -59 -175 -56 -173
rect -36 -175 -34 -172
rect -20 -176 -18 -172
rect 148 -177 150 -165
rect 156 -177 158 -165
rect 172 -177 174 -165
rect 188 -177 190 -165
rect 196 -169 198 -165
rect 196 -177 198 -174
rect 212 -177 214 -165
rect 229 -177 231 -165
rect 245 -177 247 -165
rect 261 -168 263 -165
rect 261 -177 263 -174
rect 49 -180 51 -177
rect 57 -180 59 -177
rect 73 -180 75 -177
rect 89 -180 91 -177
rect 97 -180 99 -177
rect -91 -199 -88 -197
rect -48 -199 -40 -197
rect -35 -199 -30 -197
rect 10 -199 13 -197
rect 245 -184 247 -181
rect 261 -185 263 -181
rect 172 -190 174 -187
rect 188 -190 190 -187
rect 196 -190 198 -187
rect 212 -190 214 -187
rect 229 -190 231 -187
rect 148 -200 150 -197
rect 156 -199 158 -197
rect -91 -207 -88 -205
rect -48 -207 -30 -205
rect 10 -207 13 -205
rect 49 -212 51 -200
rect 57 -212 59 -200
rect 73 -212 75 -200
rect 89 -212 91 -200
rect 97 -212 99 -200
rect -128 -226 -125 -224
rect -45 -226 -33 -224
rect 7 -226 10 -224
rect 49 -225 51 -222
rect 57 -225 59 -222
rect 73 -225 75 -222
rect -128 -234 -125 -232
rect -45 -234 -41 -232
rect -36 -234 -33 -232
rect 7 -234 10 -232
rect 89 -235 91 -232
rect 97 -234 99 -232
rect -36 -257 -34 -254
rect -20 -257 -18 -256
rect 51 -259 54 -257
rect 64 -259 67 -257
rect 148 -254 150 -251
rect 156 -254 158 -251
rect 172 -254 174 -251
rect 188 -254 190 -251
rect 196 -254 198 -251
rect 212 -254 214 -251
rect 229 -254 231 -251
rect 72 -259 76 -257
rect 96 -259 99 -257
rect -36 -269 -34 -265
rect -20 -268 -18 -265
rect 51 -267 54 -265
rect 64 -267 76 -265
rect 96 -267 99 -265
rect -35 -274 -34 -269
rect 245 -266 247 -263
rect 261 -266 263 -265
rect -36 -277 -34 -274
rect -20 -277 -18 -274
rect -104 -284 -101 -282
rect -81 -284 -69 -282
rect -59 -284 -56 -282
rect -36 -284 -34 -281
rect -20 -285 -18 -281
rect 148 -286 150 -274
rect 156 -286 158 -274
rect 172 -286 174 -274
rect 188 -286 190 -274
rect 196 -278 198 -274
rect 196 -286 198 -283
rect 212 -286 214 -274
rect 229 -286 231 -274
rect 245 -286 247 -274
rect 261 -277 263 -274
rect 261 -286 263 -283
rect 49 -289 51 -286
rect 57 -289 59 -286
rect 73 -289 75 -286
rect 89 -289 91 -286
rect 97 -289 99 -286
rect -91 -308 -88 -306
rect -48 -308 -40 -306
rect -35 -308 -30 -306
rect 10 -308 13 -306
rect 245 -293 247 -290
rect 261 -294 263 -290
rect 172 -299 174 -296
rect 188 -299 190 -296
rect 196 -299 198 -296
rect 212 -299 214 -296
rect 229 -299 231 -296
rect 148 -309 150 -306
rect 156 -308 158 -306
rect -91 -316 -88 -314
rect -48 -316 -30 -314
rect 10 -316 13 -314
rect 49 -321 51 -309
rect 57 -321 59 -309
rect 73 -321 75 -309
rect 89 -321 91 -309
rect 97 -321 99 -309
rect -128 -335 -125 -333
rect -45 -335 -33 -333
rect 7 -335 10 -333
rect 49 -334 51 -331
rect 57 -334 59 -331
rect 73 -334 75 -331
rect -128 -343 -125 -341
rect -45 -343 -41 -341
rect -36 -343 -33 -341
rect 7 -343 10 -341
rect 89 -344 91 -341
rect 97 -343 99 -341
rect -36 -366 -34 -363
rect -20 -366 -18 -365
rect 51 -368 54 -366
rect 64 -368 67 -366
rect 148 -363 150 -360
rect 156 -363 158 -360
rect 172 -363 174 -360
rect 196 -363 198 -360
rect 204 -363 206 -360
rect 72 -368 76 -366
rect 96 -368 99 -366
rect -36 -378 -34 -374
rect -20 -377 -18 -374
rect 51 -376 54 -374
rect 64 -376 76 -374
rect 96 -376 99 -374
rect -35 -383 -34 -378
rect -36 -386 -34 -383
rect -20 -386 -18 -383
rect -104 -393 -101 -391
rect -81 -393 -69 -391
rect -59 -393 -56 -391
rect -36 -393 -34 -390
rect -20 -394 -18 -390
rect 148 -395 150 -383
rect 156 -395 158 -383
rect 172 -395 174 -383
rect 49 -398 51 -395
rect 57 -398 59 -395
rect 73 -398 75 -395
rect 89 -398 91 -395
rect 97 -398 99 -395
rect -91 -417 -88 -415
rect -48 -417 -40 -415
rect -35 -417 -30 -415
rect 10 -417 13 -415
rect 216 -386 219 -384
rect 239 -386 249 -384
rect 253 -386 257 -384
rect 277 -386 280 -384
rect 216 -394 219 -392
rect 239 -394 257 -392
rect 277 -394 280 -392
rect 172 -408 174 -405
rect 196 -415 198 -403
rect 204 -407 206 -403
rect 204 -415 206 -412
rect 148 -418 150 -415
rect 156 -417 158 -415
rect -91 -425 -88 -423
rect -48 -425 -30 -423
rect 10 -425 13 -423
rect 49 -430 51 -418
rect 57 -430 59 -418
rect 73 -430 75 -418
rect 89 -430 91 -418
rect 97 -430 99 -418
rect -128 -444 -125 -442
rect -45 -444 -33 -442
rect 7 -444 10 -442
rect 49 -443 51 -440
rect 57 -443 59 -440
rect 73 -443 75 -440
rect 220 -430 223 -428
rect 243 -430 255 -428
rect 265 -430 268 -428
rect 115 -438 118 -436
rect 138 -438 156 -436
rect 176 -438 179 -436
rect 196 -438 198 -435
rect 204 -438 206 -435
rect 115 -446 118 -444
rect 138 -446 148 -444
rect 152 -446 156 -444
rect 176 -446 179 -444
rect -128 -452 -125 -450
rect -45 -452 -41 -450
rect -36 -452 -33 -450
rect 7 -452 10 -450
rect 89 -453 91 -450
rect 97 -452 99 -450
rect 192 -454 195 -452
rect 235 -454 239 -452
rect 244 -454 247 -452
rect 267 -454 270 -452
rect 192 -462 195 -460
rect 235 -462 247 -460
rect 267 -462 270 -460
<< polycontact >>
rect -22 -38 -18 -34
rect 112 -28 116 -24
rect 78 -48 82 -44
rect -124 -68 -120 -64
rect -74 -70 -70 -66
rect -22 -71 -18 -67
rect 112 -61 116 -57
rect 172 -78 176 -74
rect 45 -96 49 -92
rect -44 -102 -40 -98
rect 69 -102 73 -98
rect 85 -101 89 -97
rect -44 -115 -40 -111
rect 130 -113 134 -109
rect 172 -111 176 -107
rect 95 -129 99 -125
rect -22 -147 -18 -143
rect 71 -162 75 -158
rect 259 -156 263 -152
rect -74 -179 -70 -175
rect 144 -170 148 -166
rect -22 -180 -18 -176
rect 168 -170 172 -166
rect 184 -170 188 -166
rect 208 -176 212 -172
rect 225 -176 229 -172
rect 259 -189 263 -185
rect 45 -205 49 -201
rect -44 -211 -40 -207
rect 69 -211 73 -207
rect 85 -210 89 -206
rect 154 -203 158 -199
rect -44 -224 -40 -220
rect 95 -238 99 -234
rect -22 -256 -18 -252
rect 71 -271 75 -267
rect 259 -265 263 -261
rect -74 -288 -70 -284
rect 144 -279 148 -275
rect -22 -289 -18 -285
rect 168 -279 172 -275
rect 184 -279 188 -275
rect 208 -285 212 -281
rect 225 -285 229 -281
rect 259 -298 263 -294
rect 45 -314 49 -310
rect -44 -320 -40 -316
rect 69 -320 73 -316
rect 85 -319 89 -315
rect 154 -312 158 -308
rect -44 -333 -40 -329
rect 95 -347 99 -343
rect -22 -365 -18 -361
rect 71 -380 75 -376
rect -74 -397 -70 -393
rect 144 -388 148 -384
rect -22 -398 -18 -394
rect 168 -388 172 -384
rect 249 -387 253 -383
rect 242 -398 246 -394
rect 192 -408 196 -404
rect 45 -423 49 -419
rect -44 -429 -40 -425
rect 69 -429 73 -425
rect 85 -428 89 -424
rect 154 -421 158 -417
rect -44 -442 -40 -438
rect 141 -436 145 -432
rect 250 -434 254 -430
rect 148 -446 152 -442
rect 95 -456 99 -452
<< metal1 >>
rect 17 -22 41 -20
rect -131 -23 54 -22
rect -131 -25 20 -23
rect 38 -25 54 -23
rect 62 -21 77 -18
rect -131 -64 -128 -25
rect -125 -31 27 -28
rect 62 -28 65 -21
rect 32 -31 65 -28
rect 78 -27 112 -24
rect -125 -37 -122 -31
rect -116 -37 -109 -34
rect -116 -53 -113 -37
rect -131 -67 -124 -64
rect -116 -69 -113 -57
rect -100 -67 -97 -31
rect -46 -38 -22 -35
rect 78 -36 81 -27
rect 93 -33 96 -27
rect -46 -43 -43 -38
rect 22 -39 81 -36
rect -125 -82 -122 -79
rect -116 -93 -113 -73
rect -124 -96 -113 -93
rect -100 -91 -97 -71
rect -91 -46 -41 -43
rect -91 -77 -88 -46
rect -32 -54 -29 -47
rect -25 -52 -22 -47
rect 22 -52 25 -39
rect 78 -44 81 -39
rect 86 -49 89 -37
rect 102 -44 105 -37
rect 109 -42 112 -37
rect 109 -44 126 -42
rect 102 -45 126 -44
rect 102 -47 112 -45
rect 102 -49 105 -47
rect -25 -54 25 -52
rect -32 -55 25 -54
rect 40 -54 44 -51
rect 48 -54 70 -51
rect 89 -53 93 -50
rect 109 -49 112 -47
rect -32 -57 -22 -55
rect -32 -59 -29 -57
rect -81 -62 -69 -59
rect -65 -62 -41 -59
rect -25 -59 -22 -57
rect -41 -67 -38 -63
rect 67 -65 70 -54
rect 93 -57 96 -53
rect 93 -60 112 -57
rect -74 -77 -71 -70
rect -41 -70 -22 -67
rect 67 -68 123 -65
rect 68 -71 71 -68
rect 84 -71 87 -68
rect 101 -71 104 -68
rect -62 -74 -59 -71
rect -62 -77 14 -74
rect 120 -73 123 -68
rect 120 -76 132 -73
rect -91 -80 -68 -77
rect -88 -91 -85 -87
rect -100 -94 -85 -91
rect -100 -103 -97 -94
rect -88 -99 -85 -94
rect -132 -106 -97 -103
rect -132 -110 -129 -106
rect -71 -107 -68 -80
rect -46 -83 -27 -80
rect -46 -91 -43 -83
rect -26 -86 -16 -83
rect -48 -94 -43 -91
rect -44 -107 -41 -102
rect -71 -110 -41 -107
rect -132 -113 -125 -110
rect -132 -212 -129 -113
rect -44 -111 -41 -110
rect -33 -126 -30 -114
rect -19 -126 -16 -86
rect 11 -99 14 -77
rect 129 -82 132 -76
rect 148 -78 172 -75
rect 148 -83 151 -78
rect 148 -87 153 -83
rect 148 -89 151 -87
rect 25 -95 45 -92
rect 10 -103 14 -99
rect 61 -98 64 -91
rect 77 -98 80 -91
rect 93 -93 96 -91
rect 123 -92 151 -89
rect 123 -93 127 -92
rect 93 -96 127 -93
rect 162 -94 165 -87
rect 169 -92 172 -87
rect 169 -94 198 -92
rect 162 -95 198 -94
rect 61 -101 69 -98
rect 61 -103 64 -101
rect 77 -101 85 -98
rect 77 -103 80 -101
rect 101 -103 104 -96
rect 11 -118 14 -103
rect 48 -106 60 -103
rect 61 -112 64 -107
rect 124 -109 127 -96
rect 162 -97 172 -95
rect 162 -99 165 -97
rect 138 -107 141 -102
rect 169 -99 172 -97
rect 153 -107 156 -103
rect 124 -112 130 -109
rect 138 -110 172 -107
rect 7 -122 10 -119
rect 68 -119 71 -113
rect 138 -114 141 -110
rect 84 -119 112 -116
rect 15 -122 52 -119
rect 56 -122 84 -119
rect 117 -119 128 -116
rect 125 -120 128 -119
rect 125 -123 129 -120
rect -48 -132 -45 -130
rect -19 -129 95 -126
rect -33 -132 -29 -130
rect -48 -135 20 -132
rect 43 -137 46 -129
rect 120 -133 124 -131
rect 50 -136 124 -133
rect -46 -147 -22 -144
rect 50 -145 53 -136
rect 61 -142 80 -139
rect 61 -143 64 -142
rect -46 -152 -43 -147
rect 4 -148 53 -145
rect 76 -143 80 -142
rect -91 -155 -41 -152
rect -100 -200 -97 -180
rect -91 -186 -88 -155
rect -32 -163 -29 -156
rect -25 -161 -22 -156
rect 4 -161 7 -148
rect 15 -154 54 -151
rect -25 -163 7 -161
rect -32 -164 7 -163
rect -32 -166 -22 -164
rect -32 -168 -29 -166
rect -81 -171 -69 -168
rect -65 -171 -41 -168
rect -25 -168 -22 -166
rect -41 -176 -38 -172
rect -74 -186 -71 -179
rect -41 -179 -22 -176
rect -62 -183 -59 -180
rect 11 -183 14 -156
rect 61 -159 64 -147
rect 117 -142 227 -139
rect 80 -147 103 -144
rect 100 -154 103 -147
rect 143 -145 146 -142
rect 160 -145 163 -142
rect 167 -145 170 -142
rect 183 -145 186 -142
rect 207 -145 210 -142
rect 224 -145 227 -142
rect 100 -157 120 -154
rect 72 -166 75 -162
rect 96 -163 103 -160
rect -62 -186 14 -183
rect -91 -189 -68 -186
rect -88 -200 -85 -196
rect -100 -203 -85 -200
rect -100 -212 -97 -203
rect -88 -208 -85 -203
rect -132 -215 -97 -212
rect -132 -219 -129 -215
rect -71 -216 -68 -189
rect -46 -192 -27 -189
rect -46 -200 -43 -192
rect -26 -195 -16 -192
rect -48 -203 -43 -200
rect -44 -216 -41 -211
rect -71 -219 -41 -216
rect -132 -222 -125 -219
rect -132 -321 -129 -222
rect -44 -220 -41 -219
rect -33 -235 -30 -223
rect -19 -235 -16 -195
rect 11 -208 14 -186
rect 21 -169 75 -166
rect 21 -200 24 -169
rect 100 -180 103 -163
rect 37 -183 44 -180
rect 48 -183 68 -180
rect 72 -183 84 -180
rect 88 -183 100 -180
rect 64 -200 68 -197
rect 25 -204 45 -201
rect 10 -212 14 -208
rect 65 -207 68 -200
rect 77 -207 80 -200
rect 93 -202 96 -200
rect 117 -200 120 -157
rect 225 -155 259 -152
rect 203 -165 207 -162
rect 124 -170 144 -167
rect 152 -167 155 -165
rect 152 -170 168 -167
rect 176 -167 179 -165
rect 176 -170 184 -167
rect 160 -177 163 -170
rect 176 -177 179 -170
rect 204 -172 207 -165
rect 216 -172 219 -165
rect 225 -172 228 -155
rect 240 -161 243 -155
rect 204 -176 208 -172
rect 216 -175 225 -172
rect 204 -177 207 -176
rect 216 -177 219 -175
rect 233 -177 236 -165
rect 249 -172 252 -165
rect 256 -170 259 -165
rect 256 -172 273 -170
rect 249 -173 273 -172
rect 249 -175 259 -173
rect 249 -177 252 -175
rect 187 -180 199 -177
rect 203 -180 207 -177
rect 236 -181 240 -178
rect 256 -177 259 -175
rect 167 -190 170 -187
rect 192 -190 195 -187
rect 240 -185 243 -181
rect 207 -190 210 -187
rect 224 -190 227 -187
rect 240 -188 259 -185
rect 143 -193 227 -190
rect 93 -205 109 -202
rect 65 -211 69 -207
rect 77 -210 85 -207
rect 65 -212 68 -211
rect 77 -212 80 -210
rect 101 -212 104 -205
rect 117 -203 154 -200
rect 11 -225 14 -212
rect 48 -215 60 -212
rect 64 -215 68 -212
rect 138 -214 141 -203
rect 53 -225 56 -222
rect 68 -225 71 -222
rect 163 -225 166 -193
rect 11 -227 166 -225
rect 7 -231 10 -228
rect 15 -228 166 -227
rect -48 -241 -45 -239
rect -19 -238 95 -235
rect -33 -241 -29 -239
rect -48 -244 20 -241
rect 43 -246 46 -238
rect 120 -242 124 -239
rect 50 -245 124 -242
rect -46 -256 -22 -253
rect 50 -254 53 -245
rect 61 -251 79 -248
rect 61 -252 64 -251
rect -46 -261 -43 -256
rect 4 -257 53 -254
rect 76 -252 79 -251
rect -91 -264 -41 -261
rect -100 -309 -97 -289
rect -91 -295 -88 -264
rect -32 -272 -29 -265
rect -25 -270 -22 -265
rect 4 -270 7 -257
rect 15 -263 54 -260
rect -25 -272 7 -270
rect -32 -273 7 -272
rect -32 -275 -22 -273
rect -32 -277 -29 -275
rect -81 -280 -69 -277
rect -65 -280 -41 -277
rect -25 -277 -22 -275
rect -41 -285 -38 -281
rect -74 -295 -71 -288
rect -41 -288 -22 -285
rect -62 -292 -59 -289
rect 11 -292 14 -265
rect 61 -268 64 -256
rect 80 -255 109 -252
rect 117 -251 227 -248
rect 72 -275 75 -271
rect 96 -272 103 -269
rect -62 -295 14 -292
rect -91 -298 -68 -295
rect -88 -309 -85 -305
rect -100 -312 -85 -309
rect -100 -321 -97 -312
rect -88 -317 -85 -312
rect -132 -324 -97 -321
rect -132 -328 -129 -324
rect -71 -325 -68 -298
rect -46 -301 -27 -298
rect -46 -309 -43 -301
rect -26 -304 -16 -301
rect -48 -312 -43 -309
rect -44 -325 -41 -320
rect -71 -328 -41 -325
rect -132 -331 -125 -328
rect -132 -430 -129 -331
rect -44 -329 -41 -328
rect -33 -344 -30 -332
rect -19 -344 -16 -304
rect 11 -317 14 -295
rect 21 -278 75 -275
rect 21 -309 24 -278
rect 100 -289 103 -272
rect 106 -283 109 -255
rect 143 -254 146 -251
rect 160 -254 163 -251
rect 167 -254 170 -251
rect 183 -254 186 -251
rect 207 -254 210 -251
rect 224 -254 227 -251
rect 225 -264 259 -261
rect 203 -274 207 -271
rect 122 -279 144 -276
rect 152 -276 155 -274
rect 152 -279 168 -276
rect 176 -276 179 -274
rect 176 -279 184 -276
rect 106 -286 120 -283
rect 160 -286 163 -279
rect 176 -286 179 -279
rect 204 -281 207 -274
rect 216 -281 219 -274
rect 225 -281 228 -264
rect 240 -270 243 -264
rect 204 -285 208 -281
rect 216 -284 225 -281
rect 204 -286 207 -285
rect 216 -286 219 -284
rect 233 -286 236 -274
rect 249 -281 252 -274
rect 256 -279 259 -274
rect 256 -281 273 -279
rect 249 -282 273 -281
rect 249 -284 259 -282
rect 249 -286 252 -284
rect 37 -292 44 -289
rect 48 -292 68 -289
rect 72 -292 84 -289
rect 88 -292 100 -289
rect 64 -309 68 -306
rect 25 -313 45 -310
rect 10 -321 14 -317
rect 65 -316 68 -309
rect 77 -316 80 -309
rect 93 -311 96 -309
rect 117 -309 120 -286
rect 187 -289 199 -286
rect 203 -289 207 -286
rect 236 -290 240 -287
rect 256 -286 259 -284
rect 167 -299 170 -296
rect 192 -299 195 -296
rect 240 -294 243 -290
rect 207 -299 210 -296
rect 224 -299 227 -296
rect 240 -297 259 -294
rect 143 -302 227 -299
rect 93 -314 109 -311
rect 65 -320 69 -316
rect 77 -319 85 -316
rect 65 -321 68 -320
rect 77 -321 80 -319
rect 101 -321 104 -314
rect 117 -312 154 -309
rect 11 -334 14 -321
rect 48 -324 60 -321
rect 64 -324 68 -321
rect 53 -334 56 -331
rect 68 -334 71 -331
rect 163 -334 166 -302
rect 11 -336 166 -334
rect 7 -340 10 -337
rect 15 -337 166 -336
rect -48 -350 -45 -348
rect -19 -347 95 -344
rect -33 -350 -29 -348
rect -48 -353 20 -350
rect 43 -355 46 -347
rect 121 -351 124 -348
rect 50 -354 124 -351
rect -46 -365 -22 -362
rect 50 -363 53 -354
rect 61 -360 80 -357
rect 61 -361 64 -360
rect -46 -370 -43 -365
rect 4 -366 53 -363
rect 76 -361 80 -360
rect -91 -373 -41 -370
rect -100 -418 -97 -398
rect -91 -404 -88 -373
rect -32 -381 -29 -374
rect -25 -379 -22 -374
rect 4 -379 7 -366
rect 15 -373 54 -370
rect -25 -381 7 -379
rect -32 -382 7 -381
rect -32 -384 -22 -382
rect -32 -386 -29 -384
rect -81 -389 -69 -386
rect -65 -389 -41 -386
rect -25 -386 -22 -384
rect -41 -394 -38 -390
rect -74 -404 -71 -397
rect -41 -397 -22 -394
rect -62 -401 -59 -398
rect 11 -401 14 -374
rect 61 -377 64 -365
rect 80 -364 109 -361
rect 117 -360 215 -357
rect 72 -384 75 -380
rect 96 -381 103 -378
rect -62 -404 14 -401
rect -91 -407 -68 -404
rect -88 -418 -85 -414
rect -100 -421 -85 -418
rect -100 -430 -97 -421
rect -88 -426 -85 -421
rect -132 -433 -97 -430
rect -132 -437 -129 -433
rect -71 -434 -68 -407
rect -46 -410 -27 -407
rect -46 -418 -43 -410
rect -26 -413 -16 -410
rect -48 -421 -43 -418
rect -44 -434 -41 -429
rect -71 -437 -41 -434
rect -132 -440 -125 -437
rect -132 -463 -129 -440
rect -44 -438 -41 -437
rect -33 -453 -30 -441
rect -19 -453 -16 -413
rect 11 -426 14 -404
rect 21 -387 75 -384
rect 21 -418 24 -387
rect 100 -398 103 -381
rect 106 -392 109 -364
rect 143 -363 146 -360
rect 160 -363 163 -360
rect 167 -363 170 -360
rect 191 -363 194 -360
rect 212 -379 215 -360
rect 241 -376 244 -369
rect 241 -379 260 -376
rect 130 -385 133 -380
rect 212 -382 219 -379
rect 130 -388 144 -385
rect 152 -385 155 -383
rect 152 -388 168 -385
rect 176 -385 179 -383
rect 176 -388 190 -385
rect 106 -395 120 -392
rect 160 -395 163 -388
rect 176 -395 179 -388
rect 37 -401 44 -398
rect 48 -401 68 -398
rect 72 -401 84 -398
rect 88 -401 100 -398
rect 64 -418 68 -415
rect 25 -422 45 -419
rect 10 -430 14 -426
rect 65 -425 68 -418
rect 77 -425 80 -418
rect 93 -420 96 -418
rect 117 -418 120 -395
rect 187 -404 190 -388
rect 219 -395 222 -383
rect 241 -387 244 -379
rect 239 -390 244 -387
rect 211 -402 215 -400
rect 243 -402 246 -398
rect 211 -403 246 -402
rect 167 -408 170 -405
rect 187 -407 192 -404
rect 212 -405 246 -403
rect 143 -411 175 -408
rect 93 -423 109 -420
rect 65 -429 69 -425
rect 77 -428 85 -425
rect 65 -430 68 -429
rect 77 -430 80 -428
rect 101 -430 104 -423
rect 117 -421 154 -418
rect 11 -443 14 -430
rect 48 -433 60 -430
rect 64 -433 68 -430
rect 111 -434 118 -431
rect 53 -443 56 -440
rect 68 -443 71 -440
rect 11 -445 87 -443
rect 7 -449 11 -446
rect 16 -446 87 -445
rect 111 -448 114 -434
rect 142 -432 145 -425
rect 138 -443 143 -440
rect 111 -451 118 -448
rect 140 -451 143 -443
rect 148 -442 151 -421
rect 172 -431 175 -411
rect 212 -415 215 -405
rect 195 -418 207 -415
rect 211 -418 215 -415
rect 249 -423 252 -387
rect 263 -399 273 -396
rect 243 -426 255 -423
rect 176 -434 199 -431
rect 214 -435 223 -432
rect 263 -431 266 -399
rect -48 -459 -45 -457
rect -19 -456 95 -453
rect 111 -454 114 -451
rect 140 -454 163 -451
rect -33 -459 -29 -457
rect -48 -462 20 -459
rect 172 -467 175 -435
rect 214 -463 217 -435
rect 250 -443 253 -434
rect 265 -435 266 -431
rect 232 -446 253 -443
rect 232 -447 235 -446
rect 247 -447 251 -446
rect 183 -464 195 -463
rect 180 -466 195 -464
rect 199 -466 217 -463
rect 247 -463 250 -451
rect 263 -455 266 -435
rect 16 -470 175 -467
rect 263 -470 266 -459
rect 172 -473 266 -470
<< m2contact >>
rect 54 -25 59 -20
rect -109 -39 -104 -34
rect -126 -87 -121 -82
rect -129 -97 -124 -92
rect 20 -96 25 -91
rect 10 -123 15 -118
rect 112 -120 117 -115
rect 20 -137 25 -132
rect 120 -131 125 -126
rect 42 -142 47 -137
rect 10 -156 15 -151
rect 20 -205 25 -200
rect 123 -167 128 -162
rect 109 -206 114 -201
rect 10 -232 15 -227
rect 20 -246 25 -241
rect 120 -239 125 -234
rect 42 -251 47 -246
rect 10 -265 15 -260
rect 20 -314 25 -309
rect 109 -315 114 -310
rect 10 -341 15 -336
rect 20 -355 25 -350
rect 120 -348 125 -343
rect 42 -360 47 -355
rect 10 -374 15 -369
rect 20 -423 25 -418
rect 109 -424 114 -419
rect 11 -450 16 -445
rect 163 -455 168 -450
rect 20 -464 25 -459
rect 11 -470 16 -465
<< pm12contact >>
rect -40 -56 -35 -51
rect 56 -47 61 -42
rect 93 -45 98 -40
rect -40 -92 -35 -87
rect -41 -128 -36 -123
rect 154 -96 159 -91
rect -40 -165 -35 -160
rect 67 -150 72 -145
rect -40 -201 -35 -196
rect -41 -237 -36 -232
rect 56 -177 61 -172
rect 196 -174 201 -169
rect 240 -173 245 -168
rect -40 -274 -35 -269
rect 67 -259 72 -254
rect -40 -310 -35 -305
rect -41 -346 -36 -341
rect 56 -286 61 -281
rect 196 -283 201 -278
rect 240 -282 245 -277
rect -40 -383 -35 -378
rect 67 -368 72 -363
rect -40 -419 -35 -414
rect -41 -455 -36 -450
rect 56 -395 61 -390
rect 204 -412 209 -407
rect 239 -454 244 -449
rect 236 -467 241 -462
<< pdm12contact >>
rect -17 -47 -12 -42
rect 117 -37 122 -32
rect 177 -87 182 -82
rect -17 -156 -12 -151
rect 264 -165 269 -160
rect -17 -265 -12 -260
rect 264 -274 269 -269
rect -17 -374 -12 -369
<< ndm12contact >>
rect -17 -64 -12 -59
rect 76 -59 81 -54
rect 117 -54 122 -49
rect 177 -104 182 -99
rect -17 -173 -12 -168
rect 264 -182 269 -177
rect -17 -282 -12 -277
rect 264 -291 269 -286
rect -17 -391 -12 -386
<< metal2 >>
rect 59 -25 69 -22
rect 66 -26 69 -25
rect 66 -29 76 -26
rect -104 -38 60 -35
rect 57 -42 60 -38
rect -16 -51 -13 -47
rect -35 -54 -13 -51
rect -121 -86 -106 -83
rect -128 -474 -125 -97
rect -109 -137 -106 -86
rect -39 -87 -36 -56
rect -16 -59 -13 -54
rect -39 -123 -36 -92
rect 11 -137 14 -123
rect 21 -132 24 -96
rect 66 -123 69 -29
rect 73 -40 76 -29
rect 73 -43 93 -40
rect 118 -41 121 -37
rect 98 -44 121 -41
rect 118 -49 121 -44
rect 77 -63 80 -59
rect 77 -66 116 -63
rect 113 -115 116 -66
rect 178 -91 181 -87
rect 121 -96 154 -93
rect 159 -94 181 -91
rect 66 -126 108 -123
rect 121 -126 124 -96
rect 178 -99 181 -94
rect 34 -132 71 -130
rect 25 -133 71 -132
rect 25 -135 37 -133
rect -109 -140 14 -137
rect 11 -151 14 -140
rect -16 -160 -13 -156
rect -35 -163 -13 -160
rect -39 -196 -36 -165
rect -16 -168 -13 -163
rect 43 -172 46 -142
rect 68 -145 71 -133
rect 105 -162 108 -126
rect 105 -165 123 -162
rect 43 -175 56 -172
rect 110 -174 196 -171
rect 220 -171 240 -168
rect -39 -232 -36 -201
rect 110 -201 113 -174
rect 130 -178 133 -174
rect 11 -260 14 -232
rect 21 -241 24 -205
rect 220 -207 223 -171
rect 265 -169 268 -165
rect 245 -172 268 -169
rect 265 -177 268 -172
rect 121 -210 223 -207
rect 121 -234 124 -210
rect 35 -241 71 -239
rect 25 -242 71 -241
rect 25 -244 38 -242
rect -16 -269 -13 -265
rect -35 -272 -13 -269
rect -39 -305 -36 -274
rect -16 -277 -13 -272
rect 43 -281 46 -251
rect 68 -254 71 -242
rect 43 -284 56 -281
rect 110 -283 196 -280
rect 220 -280 240 -277
rect -39 -341 -36 -310
rect 110 -310 113 -283
rect 11 -369 14 -341
rect 21 -350 24 -314
rect 220 -316 223 -280
rect 265 -278 268 -274
rect 245 -281 268 -278
rect 265 -286 268 -281
rect 121 -319 223 -316
rect 121 -343 124 -319
rect 35 -350 71 -348
rect 25 -351 71 -350
rect 25 -353 38 -351
rect -16 -378 -13 -374
rect -35 -381 -13 -378
rect -39 -414 -36 -383
rect -16 -386 -13 -381
rect 43 -391 46 -360
rect 68 -363 71 -351
rect 43 -394 56 -391
rect 110 -392 186 -389
rect -39 -450 -36 -419
rect 110 -419 113 -392
rect 183 -409 186 -392
rect 183 -412 204 -409
rect 11 -465 14 -450
rect 21 -459 24 -423
rect 168 -454 190 -451
rect 187 -455 190 -454
rect 239 -455 242 -454
rect 187 -458 242 -455
rect 237 -474 240 -467
rect -128 -477 240 -474
<< m123contact >>
rect 27 -31 32 -26
rect 35 -55 40 -50
rect 121 -89 126 -84
rect 112 -144 117 -139
rect 32 -185 37 -180
rect 129 -183 134 -178
rect 137 -219 142 -214
rect 112 -253 117 -248
rect 121 -276 126 -271
rect 32 -293 37 -288
rect 112 -362 117 -357
rect 129 -380 134 -375
rect 32 -402 37 -397
rect 137 -429 142 -424
rect 110 -459 115 -454
rect 178 -464 183 -459
<< metal3 >>
rect 28 -51 31 -31
rect 28 -54 35 -51
rect 28 -139 31 -54
rect 28 -142 112 -139
rect 28 -180 31 -142
rect 28 -185 32 -180
rect 28 -248 31 -185
rect 28 -251 112 -248
rect 28 -288 31 -251
rect 122 -271 125 -89
rect 28 -293 32 -288
rect 28 -357 31 -293
rect 28 -360 112 -357
rect 28 -397 31 -360
rect 130 -375 133 -183
rect 28 -402 32 -397
rect 28 -459 31 -402
rect 138 -424 141 -219
rect 28 -462 178 -459
<< labels >>
rlabel metal1 17 -243 17 -243 1 Pt1
rlabel metal1 17 -352 17 -352 1 Pt2
rlabel metal1 18 -461 18 -461 1 Pt3
rlabel metal1 18 -455 18 -455 1 G3
rlabel metal1 17 -346 17 -346 1 G2
rlabel metal1 17 -237 17 -237 1 G1
rlabel metal2 -37 -436 -37 -436 1 B_3
rlabel metal1 -43 -436 -43 -436 1 A_3
rlabel metal2 -38 -327 -38 -327 1 B_2
rlabel metal1 -42 -327 -42 -327 1 A_2
rlabel metal2 -38 -217 -38 -217 1 B_1
rlabel metal1 -42 -217 -42 -217 1 A_1
rlabel metal1 -131 -443 -131 -443 3 VDD
rlabel metal1 13 -332 13 -332 7 gnd
rlabel metal1 -131 -334 -131 -334 3 VDD
rlabel metal1 16 -54 16 -54 1 pgxor0
rlabel metal1 13 -114 13 -114 7 gnd
rlabel metal1 -131 -116 -131 -116 3 VDD
rlabel metal1 13 -223 13 -223 7 gnd
rlabel metal1 -131 -225 -131 -225 3 VDD
rlabel metal1 -43 -109 -43 -109 1 A_0
rlabel metal2 -38 -109 -38 -109 1 B_0
rlabel metal1 17 -134 17 -134 1 Pt0
rlabel metal1 17 -128 17 -128 1 G0
rlabel metal1 39 -203 39 -203 1 Pt1
rlabel metal1 61 -227 61 -227 1 gnd
rlabel metal1 61 -336 61 -336 1 gnd
rlabel m2contact 112 -313 112 -313 7 GPG2
rlabel metal1 39 -312 39 -312 1 Pt2
rlabel metal1 39 -421 39 -421 1 Pt3
rlabel metal1 56 -346 56 -346 1 G2
rlabel metal2 -120 -84 -120 -84 1 gnd
rlabel metal1 -123 -29 -123 -29 5 VDD
rlabel metal1 -115 -67 -115 -67 1 C0bar
rlabel metal1 -129 -66 -129 -66 3 C0
rlabel metal2 48 -37 48 -37 1 C0bar
rlabel metal1 118 -95 118 -95 1 C1
rlabel metal2 52 -174 52 -174 1 G0
rlabel metal1 115 -135 115 -135 1 pgxor1
rlabel metal1 131 -74 131 -74 5 VDD
rlabel metal1 109 -118 109 -118 1 gnd
rlabel metal1 193 -94 193 -94 7 S1
rlabel metal1 101 -162 101 -162 1 VDD
rlabel metal1 6 -163 6 -163 1 pgxor1
rlabel metal1 64 -141 64 -141 1 P10
rlabel metal1 107 -204 107 -204 1 GPG1
rlabel metal2 126 -173 126 -173 1 GPG1
rlabel metal2 51 -283 51 -283 1 G1
rlabel metal1 4 -272 4 -272 1 pgxor2
rlabel metal1 126 -169 126 -169 1 C0
rlabel metal1 125 -202 125 -202 1 P10
rlabel metal1 114 -244 114 -244 1 pgxor2
rlabel metal2 51 -393 51 -393 1 G2
rlabel metal1 4 -381 4 -381 1 pgxor3
rlabel metal1 50 -372 50 -372 1 gnd
rlabel metal1 125 -44 125 -44 1 S0
rlabel metal2 67 -24 67 -24 1 C0
rlabel metal2 125 -282 125 -282 1 GPG2
rlabel metal1 125 -278 125 -278 1 C1
rlabel m2contact 111 -422 111 -422 7 GPG3
rlabel metal1 127 -420 127 -420 1 P32
rlabel metal3 123 -151 123 -151 1 C1
rlabel metal3 131 -295 131 -295 1 GPG1
rlabel metal1 61 -445 61 -445 1 gnd
rlabel metal1 13 -441 13 -441 7 gnd
rlabel metal1 101 -380 101 -380 1 VDD
rlabel metal2 130 -391 130 -391 1 GPG3
rlabel metal1 271 -172 271 -172 1 S2
rlabel metal2 221 -184 221 -184 1 pgxor2
rlabel metal1 187 -192 187 -192 1 gnd
rlabel metal1 149 -140 149 -140 5 VDD
rlabel metal2 222 -292 222 -292 1 pgxor3
rlabel metal1 272 -281 272 -281 1 S3
rlabel metal1 187 -301 187 -301 1 gnd
rlabel metal1 149 -249 149 -249 5 VDD
rlabel metal1 112 -437 112 -437 3 VDD
rlabel metal1 174 -438 174 -438 7 gnd
rlabel metal3 140 -330 140 -330 1 P10
rlabel metal2 179 -453 179 -453 1 Pout
rlabel metal2 179 -476 179 -476 1 C0bar
rlabel metal1 264 -471 264 -471 1 gnd
rlabel metal1 186 -465 186 -465 1 VDD
rlabel metal1 215 -433 215 -433 3 VDD
rlabel metal1 216 -404 216 -404 1 Gout
rlabel metal1 243 -371 243 -371 1 C4
rlabel metal1 265 -403 265 -403 1 gnd
rlabel metal1 208 -358 208 -358 1 VDD
rlabel metal1 131 -387 131 -387 1 GPG1
rlabel metal1 217 -283 217 -283 1 C3
rlabel metal1 218 -174 218 -174 1 C2
rlabel metal1 123 -350 123 -350 1 pgxor3
rlabel metal3 29 -183 29 -183 1 VDD
rlabel metal3 30 -291 30 -291 1 VDD
rlabel metal2 69 -253 69 -253 1 Pt1
rlabel metal1 68 -277 68 -277 1 Pt2
rlabel metal1 50 -262 50 -262 1 gnd
rlabel metal1 107 -255 107 -255 1 P21
rlabel metal1 101 -271 101 -271 1 VDD
<< end >>
