magic
tech scmos
timestamp 1731491580
<< nwell >>
rect -196 -47 -124 -15
<< ntransistor >>
rect -185 -63 -183 -53
rect -177 -63 -175 -53
rect -161 -63 -159 -53
rect -145 -73 -143 -53
rect -137 -73 -135 -53
<< ptransistor >>
rect -185 -41 -183 -21
rect -177 -41 -175 -21
rect -161 -41 -159 -21
rect -145 -41 -143 -21
rect -137 -41 -135 -21
<< ndiffusion >>
rect -186 -57 -185 -53
rect -190 -63 -185 -57
rect -183 -59 -177 -53
rect -183 -63 -182 -59
rect -178 -63 -177 -59
rect -175 -57 -174 -53
rect -175 -63 -170 -57
rect -166 -59 -161 -53
rect -162 -63 -161 -59
rect -159 -57 -158 -53
rect -159 -63 -154 -57
rect -150 -69 -145 -53
rect -146 -73 -145 -69
rect -143 -73 -137 -53
rect -135 -57 -134 -53
rect -135 -73 -130 -57
<< pdiffusion >>
rect -186 -25 -185 -21
rect -190 -41 -185 -25
rect -183 -41 -177 -21
rect -175 -37 -170 -21
rect -175 -41 -174 -37
rect -162 -25 -161 -21
rect -166 -41 -161 -25
rect -159 -37 -154 -21
rect -159 -41 -158 -37
rect -146 -25 -145 -21
rect -150 -41 -145 -25
rect -143 -37 -137 -21
rect -143 -41 -142 -37
rect -138 -41 -137 -37
rect -135 -25 -134 -21
rect -135 -41 -130 -25
<< ndcontact >>
rect -190 -57 -186 -53
rect -182 -63 -178 -59
rect -174 -57 -170 -53
rect -166 -63 -162 -59
rect -158 -57 -154 -53
rect -150 -73 -146 -69
rect -134 -57 -130 -53
<< pdcontact >>
rect -190 -25 -186 -21
rect -174 -41 -170 -37
rect -166 -25 -162 -21
rect -158 -41 -154 -37
rect -150 -25 -146 -21
rect -142 -41 -138 -37
rect -134 -25 -130 -21
<< polysilicon >>
rect -185 -21 -183 -18
rect -177 -21 -175 -18
rect -161 -21 -159 -18
rect -145 -21 -143 -18
rect -137 -21 -135 -18
rect -185 -53 -183 -41
rect -177 -45 -175 -41
rect -177 -53 -175 -50
rect -161 -53 -159 -41
rect -145 -53 -143 -41
rect -137 -53 -135 -41
rect -185 -66 -183 -63
rect -177 -66 -175 -63
rect -161 -66 -159 -63
rect -145 -76 -143 -73
rect -137 -75 -135 -73
<< polycontact >>
rect -189 -46 -185 -42
rect -165 -52 -161 -48
rect -149 -51 -145 -47
rect -139 -79 -135 -75
<< metal1 >>
rect -196 -18 -124 -15
rect -190 -21 -187 -18
rect -166 -21 -163 -18
rect -150 -21 -147 -18
rect -133 -21 -130 -18
rect -170 -41 -166 -38
rect -198 -45 -189 -42
rect -169 -48 -166 -41
rect -157 -48 -154 -41
rect -141 -43 -138 -41
rect -141 -46 -119 -43
rect -169 -52 -165 -48
rect -157 -51 -149 -48
rect -169 -53 -166 -52
rect -157 -53 -154 -51
rect -186 -56 -174 -53
rect -170 -56 -166 -53
rect -130 -56 -127 -46
rect -181 -66 -178 -63
rect -166 -66 -163 -63
rect -188 -69 -147 -66
rect -198 -79 -139 -76
<< pm12contact >>
rect -177 -50 -172 -45
<< metal2 >>
rect -198 -50 -177 -47
<< labels >>
rlabel metal1 -127 -45 -127 -45 1 out
rlabel metal1 -184 -16 -184 -16 5 VDD
rlabel metal1 -186 -68 -186 -68 1 gnd
rlabel metal1 -197 -78 -197 -78 3 interNAND
rlabel metal2 -197 -49 -197 -49 3 interORg
rlabel metal1 -197 -44 -197 -44 3 interORp
<< end >>
