magic
tech scmos
timestamp 1731450193
<< nwell >>
rect -210 143 -178 180
rect 16 173 28 176
rect -210 88 -151 143
rect 4 141 28 173
rect -125 100 -93 120
rect 44 105 64 146
rect -125 96 -90 100
rect -166 85 -151 88
rect -110 55 -90 96
<< ntransistor >>
rect 15 125 17 135
rect 34 133 38 135
rect 34 117 38 119
rect -141 107 -131 109
rect -199 42 -197 82
rect -191 42 -189 82
rect -120 83 -116 85
rect -172 39 -170 79
rect -164 39 -162 79
rect -120 67 -116 69
<< ptransistor >>
rect -199 94 -197 174
rect -191 94 -189 174
rect 15 147 17 167
rect -172 97 -170 137
rect -164 97 -162 137
rect 50 133 58 135
rect 50 117 58 119
rect -119 107 -99 109
rect -104 83 -96 85
rect -104 67 -96 69
<< ndiffusion >>
rect 34 135 38 136
rect 10 129 15 135
rect 14 125 15 129
rect 17 131 18 135
rect 17 125 22 131
rect 34 132 38 133
rect 34 119 38 120
rect 34 116 38 117
rect -137 110 -131 114
rect -141 109 -131 110
rect -141 106 -131 107
rect -141 102 -135 106
rect -200 78 -199 82
rect -204 42 -199 78
rect -197 46 -191 82
rect -197 42 -196 46
rect -192 42 -191 46
rect -189 78 -188 82
rect -120 85 -116 86
rect -120 82 -116 83
rect -189 42 -184 78
rect -177 43 -172 79
rect -173 39 -172 43
rect -170 39 -164 79
rect -162 75 -161 79
rect -162 39 -157 75
rect -120 69 -116 70
rect -120 66 -116 67
<< pdiffusion >>
rect -204 98 -199 174
rect -200 94 -199 98
rect -197 94 -191 174
rect -189 170 -188 174
rect -189 94 -184 170
rect 14 163 15 167
rect 10 147 15 163
rect 17 151 22 167
rect 17 147 18 151
rect -173 133 -172 137
rect -177 97 -172 133
rect -170 101 -164 137
rect -170 97 -169 101
rect -165 97 -164 101
rect -162 133 -161 137
rect -162 97 -157 133
rect 54 136 58 140
rect 50 135 58 136
rect 50 132 58 133
rect 54 128 58 132
rect 54 120 58 124
rect 50 119 58 120
rect -119 110 -103 114
rect 50 116 58 117
rect 55 112 58 116
rect -119 109 -99 110
rect -119 106 -99 107
rect -115 102 -99 106
rect -100 86 -96 90
rect -104 85 -96 86
rect -104 82 -96 83
rect -100 78 -96 82
rect -100 70 -96 74
rect -104 69 -96 70
rect -104 66 -96 67
rect -99 62 -96 66
<< ndcontact >>
rect 34 136 38 140
rect 10 125 14 129
rect 18 131 22 135
rect 34 128 38 132
rect 34 120 38 124
rect -141 110 -137 114
rect -135 102 -131 106
rect -204 78 -200 82
rect -196 42 -192 46
rect -188 78 -184 82
rect -120 86 -116 90
rect -177 39 -173 43
rect -161 75 -157 79
rect -120 78 -116 82
rect -120 70 -116 74
<< pdcontact >>
rect -204 94 -200 98
rect -188 170 -184 174
rect 10 163 14 167
rect 18 147 22 151
rect -177 133 -173 137
rect -169 97 -165 101
rect -161 133 -157 137
rect 50 136 54 140
rect 50 128 54 132
rect 50 120 54 124
rect -103 110 -99 114
rect -119 102 -115 106
rect -104 86 -100 90
rect -104 78 -100 82
rect -104 70 -100 74
<< polysilicon >>
rect -199 174 -197 177
rect -191 174 -189 177
rect 15 167 17 170
rect -172 137 -170 140
rect -164 137 -162 140
rect 15 135 17 147
rect 31 133 34 135
rect 38 134 41 135
rect 46 134 50 135
rect 38 133 50 134
rect 58 133 61 135
rect 15 122 17 125
rect 29 117 34 119
rect 38 117 41 119
rect 47 117 50 119
rect 58 117 59 119
rect -144 107 -141 109
rect -131 107 -119 109
rect -99 107 -96 109
rect -199 90 -197 94
rect -199 82 -197 85
rect -191 82 -189 94
rect -172 79 -170 97
rect -164 89 -162 97
rect -164 79 -162 84
rect -123 83 -120 85
rect -116 84 -113 85
rect -108 84 -104 85
rect -116 83 -104 84
rect -96 83 -93 85
rect -199 39 -197 42
rect -191 39 -189 42
rect -124 67 -120 69
rect -116 67 -113 69
rect -107 67 -104 69
rect -96 67 -95 69
rect -172 36 -170 39
rect -164 36 -162 39
<< polycontact >>
rect 11 136 15 140
rect 25 117 29 121
rect 59 117 63 121
rect -130 109 -126 113
rect -189 89 -185 93
rect -176 89 -172 93
rect -128 67 -124 71
rect -95 67 -91 71
<< metal1 >>
rect -210 178 -178 181
rect -187 174 -184 178
rect 4 173 28 176
rect 10 167 13 173
rect 5 157 54 160
rect 5 140 8 157
rect 19 142 22 147
rect 51 145 54 157
rect 51 142 62 145
rect 19 140 29 142
rect 51 140 54 142
rect 5 137 11 140
rect -173 134 -161 137
rect 19 139 34 140
rect 19 135 22 139
rect 26 137 34 139
rect 10 122 13 125
rect -184 119 -126 120
rect -184 117 -106 119
rect -208 94 -204 97
rect -208 82 -205 94
rect -184 93 -181 117
rect -129 116 -106 117
rect -147 111 -141 114
rect -147 102 -144 111
rect -129 113 -126 116
rect -131 102 -119 105
rect -168 95 -165 97
rect -185 90 -176 93
rect -168 92 -150 95
rect -208 79 -204 82
rect -200 79 -188 82
rect -157 76 -154 92
rect -127 90 -124 102
rect -109 95 -106 116
rect -93 114 -90 120
rect 10 119 22 122
rect 26 121 29 137
rect 38 128 50 131
rect 40 124 43 128
rect 38 121 50 124
rect -99 111 -90 114
rect -93 100 -90 111
rect 42 107 45 121
rect 59 121 62 142
rect -109 92 -92 95
rect -104 90 -100 92
rect -127 87 -120 90
rect -127 71 -124 87
rect -116 78 -104 81
rect -114 74 -111 78
rect -116 71 -104 74
rect -112 57 -109 71
rect -95 71 -92 92
rect -196 38 -193 42
rect -205 35 -184 38
rect -177 35 -174 39
rect -177 32 -158 35
<< pm12contact >>
rect -202 85 -197 90
rect -166 84 -161 89
rect 41 134 46 139
rect -113 84 -108 89
<< pdm12contact >>
rect 50 111 55 116
rect -104 61 -99 66
<< ndm12contact >>
rect 33 111 38 116
rect -121 61 -116 66
<< metal2 >>
rect 2 153 44 156
rect 41 139 44 153
rect 43 115 46 134
rect 38 112 50 115
rect -197 85 -166 88
rect -161 85 -113 88
rect -111 65 -108 84
rect -116 62 -104 65
use XOR  XOR_0
timestamp 1731446490
transform 1 0 274 0 1 237
box -351 -83 -274 -26
<< labels >>
rlabel metal1 -188 36 -188 36 1 gnd
rlabel metal1 -190 180 -190 180 5 VDD
rlabel metal1 -206 86 -206 86 3 out
rlabel metal1 -182 91 -182 91 7 A
rlabel metal2 -182 86 -182 86 7 B
rlabel metal1 43 108 43 108 3 out
rlabel metal1 12 175 12 175 5 VDD
rlabel metal1 15 120 15 120 1 gnd
rlabel metal1 7 138 7 138 1 A
rlabel metal1 -91 112 -91 112 7 VDD
rlabel metal1 -146 109 -146 109 3 gnd
rlabel metal1 -128 117 -128 117 3 A
rlabel metal1 -111 58 -111 58 3 out
<< end >>
