* SPICE3 file created from TSPC2.ext - technology: scmos

.option scale=0.09u

M1000 a_380_n536# clk a_380_n568# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=80 ps=48
M1001 a_380_n568# mid gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=300 ps=160
M1002 a_402_n568# a_380_n536# gnd Gnd nfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1003 a_380_n536# mid VDD w_323_n542# pfet w=20 l=2
+  ad=100 pd=50 as=600 ps=280
M1004 Q clk a_402_n568# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1005 Q a_380_n536# VDD w_323_n542# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1006 mid clk a_358_n536# w_323_n542# pfet w=40 l=2
+  ad=200 pd=90 as=160 ps=88
M1007 a_358_n536# a_336_n558# VDD w_323_n542# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_336_n558# clk a_336_n536# w_323_n542# pfet w=40 l=2
+  ad=200 pd=90 as=160 ps=88
M1009 a_336_n536# D VDD w_323_n542# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 mid a_336_n558# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1011 a_336_n558# D gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 Q w_323_n542# 0.03fF
C1 w_323_n542# mid 0.09fF
C2 w_323_n542# clk 0.45fF
C3 mid clk 0.33fF
C4 w_323_n542# D 0.06fF
C5 D clk 0.03fF
C6 w_323_n542# VDD 0.08fF
C7 mid VDD 0.08fF
C8 VDD clk 0.21fF
C9 mid gnd 0.06fF
C10 a_380_n536# w_323_n542# 0.11fF
C11 gnd clk 0.36fF
C12 a_380_n536# clk 0.09fF
C13 w_323_n542# a_336_n558# 0.09fF
C14 a_336_n558# clk 0.03fF
C15 D VDD 0.06fF
C16 D gnd 0.04fF
C17 a_380_n568# gnd 0.01fF
C18 a_380_n536# VDD 0.02fF
C19 a_358_n536# VDD 0.01fF
C20 a_380_n536# gnd 0.02fF
C21 a_336_n536# VDD 0.01fF
C22 a_336_n558# VDD 0.08fF
C23 a_336_n558# gnd 0.04fF
C24 gnd Gnd 0.16fF
C25 Q Gnd 0.05fF
C26 a_380_n536# Gnd 0.11fF
C27 mid Gnd 0.13fF
C28 VDD Gnd 0.00fF
C29 a_336_n558# Gnd 0.16fF
C30 clk Gnd 0.36fF
C31 D Gnd 0.12fF
C32 w_323_n542# Gnd 3.94fF
