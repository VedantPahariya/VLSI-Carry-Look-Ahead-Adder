magic
tech scmos
timestamp 1731675722
<< nwell >>
rect 444 -378 536 -346
rect 484 -398 536 -378
<< ntransistor >>
rect 449 -340 451 -320
rect 455 -340 457 -320
rect 473 -340 475 -320
rect 479 -340 481 -320
rect 501 -340 503 -330
rect 523 -340 525 -330
<< ptransistor >>
rect 455 -372 457 -352
rect 479 -372 481 -352
rect 495 -392 497 -352
rect 501 -392 503 -352
rect 517 -392 519 -352
rect 523 -392 525 -352
<< ndiffusion >>
rect 444 -336 449 -320
rect 448 -340 449 -336
rect 451 -340 455 -320
rect 457 -324 462 -320
rect 457 -328 458 -324
rect 457 -340 462 -328
rect 468 -336 473 -320
rect 472 -340 473 -336
rect 475 -340 479 -320
rect 481 -324 486 -320
rect 481 -328 482 -324
rect 481 -340 486 -328
rect 496 -336 501 -330
rect 500 -340 501 -336
rect 503 -334 504 -330
rect 503 -340 508 -334
rect 518 -336 523 -330
rect 522 -340 523 -336
rect 525 -334 526 -330
rect 525 -340 530 -334
<< pdiffusion >>
rect 454 -356 455 -352
rect 450 -372 455 -356
rect 457 -366 462 -352
rect 457 -370 458 -366
rect 457 -372 462 -370
rect 478 -356 479 -352
rect 474 -372 479 -356
rect 481 -366 486 -352
rect 481 -370 482 -366
rect 481 -372 486 -370
rect 494 -356 495 -352
rect 490 -392 495 -356
rect 497 -392 501 -352
rect 503 -376 508 -352
rect 503 -380 504 -376
rect 503 -392 508 -380
rect 516 -356 517 -352
rect 512 -392 517 -356
rect 519 -392 523 -352
rect 525 -376 530 -352
rect 525 -380 526 -376
rect 525 -392 530 -380
<< ndcontact >>
rect 444 -340 448 -336
rect 458 -328 462 -324
rect 468 -340 472 -336
rect 482 -328 486 -324
rect 496 -340 500 -336
rect 504 -334 508 -330
rect 518 -340 522 -336
rect 526 -334 530 -330
<< pdcontact >>
rect 450 -356 454 -352
rect 458 -370 462 -366
rect 474 -356 478 -352
rect 482 -370 486 -366
rect 490 -356 494 -352
rect 504 -380 508 -376
rect 512 -356 516 -352
rect 526 -380 530 -376
<< polysilicon >>
rect 449 -320 451 -319
rect 455 -320 457 -316
rect 473 -320 475 -319
rect 479 -320 481 -316
rect 501 -330 503 -327
rect 523 -330 525 -327
rect 449 -343 451 -340
rect 455 -352 457 -340
rect 473 -343 475 -340
rect 479 -352 481 -340
rect 495 -352 497 -349
rect 501 -352 503 -340
rect 517 -352 519 -349
rect 523 -352 525 -340
rect 455 -375 457 -372
rect 479 -375 481 -372
rect 495 -399 497 -392
rect 501 -395 503 -392
rect 517 -403 519 -392
rect 523 -393 525 -392
<< polycontact >>
rect 447 -319 451 -315
rect 471 -319 475 -315
rect 457 -345 461 -341
rect 481 -350 485 -346
rect 503 -345 507 -341
rect 494 -403 498 -399
rect 513 -403 517 -399
rect 523 -397 527 -393
<< metal1 >>
rect 451 -318 471 -315
rect 475 -318 485 -315
rect 442 -327 458 -324
rect 462 -327 482 -324
rect 486 -327 530 -324
rect 505 -330 508 -327
rect 527 -330 530 -327
rect 490 -340 496 -337
rect 512 -340 518 -337
rect 444 -346 447 -340
rect 468 -342 471 -340
rect 461 -345 471 -342
rect 444 -349 453 -346
rect 444 -360 447 -349
rect 450 -352 453 -349
rect 468 -352 471 -345
rect 490 -346 493 -340
rect 512 -342 515 -340
rect 507 -345 515 -342
rect 485 -349 493 -346
rect 490 -352 493 -349
rect 512 -352 515 -345
rect 468 -355 474 -352
rect 442 -363 549 -360
rect 442 -369 458 -366
rect 462 -369 482 -366
rect 475 -377 478 -369
rect 475 -380 504 -377
rect 508 -380 526 -377
rect 476 -396 523 -393
rect 490 -403 494 -400
rect 498 -403 513 -400
<< m2contact >>
rect 485 -320 490 -315
rect 485 -404 490 -399
<< metal2 >>
rect 487 -399 490 -320
<< labels >>
rlabel metal1 514 -325 514 -325 5 gnd
rlabel metal1 508 -401 508 -401 1 clk
rlabel metal1 544 -362 544 -362 7 Q
rlabel metal1 477 -394 477 -394 1 D
rlabel metal1 469 -368 469 -368 1 VDD
<< end >>
