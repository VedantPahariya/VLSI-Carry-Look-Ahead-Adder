* SPICE3 file created from Low_Level_Latch.ext - technology: scmos

.include TSMC_180nm.txt
.option scale=0.09u
.param SUPPLY=1.8
.global gnd vdd
Vdd vdd gnd 'SUPPLY'

M1000 out clk a_14_14# w_n21_8# CMOSP w=40 l=2
+  ad=200 pd=90 as=160 ps=88
M1001 a_n8_n9# clk a_n8_14# w_n21_8# CMOSP w=40 l=2
+  ad=200 pd=90 as=160 ps=88
M1002 a_n8_14# D VDD w_n21_8# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1003 out a_n8_n9# gnd Gnd CMOSN w=11 l=2
+  ad=55 pd=32 as=110 ps=64
M1004 a_n8_n9# D gnd Gnd CMOSN w=11 l=2
+  ad=55 pd=32 as=0 ps=0
M1005 a_14_14# a_n8_n9# VDD w_n21_8# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
C0 VDD w_n21_8# 0.08fF
C1 w_n21_8# a_n8_n9# 0.09fF
C2 gnd D 0.02fF
C3 VDD clk 0.20fF
C4 w_n21_8# clk 0.13fF
C5 a_n8_n9# clk 0.03fF
C6 w_n21_8# out 0.02fF
C7 VDD D 0.05fF
C8 w_n21_8# D 0.06fF
C9 D clk 0.03fF
C10 gnd Gnd 0.09fF
C11 out Gnd 0.05fF
C12 a_n8_n9# Gnd 0.16fF
C13 clk Gnd 0.14fF
C14 D Gnd 0.12fF
C15 w_n21_8# Gnd 2.72fF

.tran 0.1n 20n
V1 clk gnd PULSE 0 'SUPPLY' 0 50p 50p 1n 2n
V2 D gnd PULSE 0 'SUPPLY' 0 50p 50p 1.75n 3.5n

.control
run
plot V(out) V(clk)+3 V(D)+6
.endc
