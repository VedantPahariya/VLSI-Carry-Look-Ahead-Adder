magic
tech scmos
timestamp 1731669992
<< nwell >>
rect 330 -548 420 -516
rect 368 -568 420 -548
<< ntransistor >>
rect 335 -510 337 -490
rect 341 -510 343 -490
rect 357 -510 359 -490
rect 363 -510 365 -490
rect 385 -510 387 -500
rect 407 -510 409 -500
<< ptransistor >>
rect 341 -542 343 -522
rect 363 -542 365 -522
rect 379 -562 381 -522
rect 385 -562 387 -522
rect 401 -562 403 -522
rect 407 -562 409 -522
<< ndiffusion >>
rect 330 -506 335 -490
rect 334 -510 335 -506
rect 337 -510 341 -490
rect 343 -494 348 -490
rect 343 -498 344 -494
rect 343 -510 348 -498
rect 352 -506 357 -490
rect 356 -510 357 -506
rect 359 -510 363 -490
rect 365 -494 370 -490
rect 365 -498 366 -494
rect 365 -510 370 -498
rect 380 -506 385 -500
rect 384 -510 385 -506
rect 387 -504 388 -500
rect 387 -510 392 -504
rect 402 -506 407 -500
rect 406 -510 407 -506
rect 409 -504 410 -500
rect 409 -510 414 -504
<< pdiffusion >>
rect 340 -526 341 -522
rect 336 -542 341 -526
rect 343 -536 348 -522
rect 343 -540 344 -536
rect 343 -542 348 -540
rect 362 -526 363 -522
rect 358 -542 363 -526
rect 365 -536 370 -522
rect 365 -540 366 -536
rect 365 -542 370 -540
rect 378 -526 379 -522
rect 374 -562 379 -526
rect 381 -562 385 -522
rect 387 -558 392 -522
rect 387 -562 388 -558
rect 400 -526 401 -522
rect 396 -562 401 -526
rect 403 -562 407 -522
rect 409 -558 414 -522
rect 409 -562 410 -558
<< ndcontact >>
rect 330 -510 334 -506
rect 344 -498 348 -494
rect 352 -510 356 -506
rect 366 -498 370 -494
rect 380 -510 384 -506
rect 388 -504 392 -500
rect 402 -510 406 -506
rect 410 -504 414 -500
<< pdcontact >>
rect 336 -526 340 -522
rect 344 -540 348 -536
rect 358 -526 362 -522
rect 366 -540 370 -536
rect 374 -526 378 -522
rect 388 -562 392 -558
rect 396 -526 400 -522
rect 410 -562 414 -558
<< polysilicon >>
rect 335 -490 337 -489
rect 341 -490 343 -486
rect 357 -490 359 -489
rect 363 -490 365 -486
rect 385 -500 387 -497
rect 407 -500 409 -497
rect 335 -513 337 -510
rect 341 -522 343 -510
rect 357 -513 359 -510
rect 363 -522 365 -510
rect 379 -522 381 -519
rect 385 -522 387 -510
rect 401 -522 403 -519
rect 407 -522 409 -510
rect 341 -545 343 -542
rect 363 -545 365 -542
rect 379 -569 381 -562
rect 385 -565 387 -562
rect 401 -573 403 -562
rect 407 -565 409 -562
<< polycontact >>
rect 333 -489 337 -485
rect 355 -489 359 -485
rect 343 -515 347 -511
rect 365 -515 369 -511
rect 387 -515 391 -511
rect 409 -515 413 -511
rect 378 -573 382 -569
rect 397 -573 401 -569
<< metal1 >>
rect 337 -488 355 -485
rect 359 -488 369 -485
rect 348 -497 366 -494
rect 370 -497 414 -494
rect 389 -500 392 -497
rect 411 -500 414 -497
rect 374 -510 380 -507
rect 396 -510 402 -507
rect 330 -512 333 -510
rect 323 -515 333 -512
rect 352 -512 355 -510
rect 347 -515 355 -512
rect 374 -512 377 -510
rect 369 -515 377 -512
rect 396 -512 399 -510
rect 391 -515 399 -512
rect 413 -515 419 -512
rect 330 -522 333 -515
rect 352 -522 355 -515
rect 374 -522 377 -515
rect 396 -522 399 -515
rect 330 -525 336 -522
rect 352 -525 358 -522
rect 348 -540 366 -537
rect 370 -540 391 -537
rect 388 -558 391 -540
rect 392 -562 410 -559
rect 375 -573 378 -570
rect 382 -573 397 -570
<< m2contact >>
rect 369 -490 374 -485
rect 370 -573 375 -568
<< metal2 >>
rect 371 -568 374 -490
<< labels >>
rlabel metal1 417 -513 417 -513 7 D
rlabel metal1 398 -495 398 -495 5 gnd
rlabel metal1 392 -571 392 -571 1 clk
rlabel metal1 324 -514 324 -514 1 Q
rlabel metal1 395 -560 395 -560 1 VDD
<< end >>
