magic
tech scmos
timestamp 1731491278
<< nwell >>
rect -77 -12 -45 20
rect -93 -74 -21 -42
rect 2 -73 90 -41
<< ntransistor >>
rect -66 -28 -64 -18
rect -58 -28 -56 -18
rect -82 -90 -80 -80
rect -74 -90 -72 -80
rect -58 -90 -56 -80
rect -42 -100 -40 -80
rect -34 -100 -32 -80
rect 13 -99 15 -79
rect 21 -99 23 -79
rect 37 -89 39 -79
rect 53 -89 55 -79
rect 61 -89 63 -79
rect 77 -89 79 -79
<< ptransistor >>
rect -66 -6 -64 14
rect -58 -6 -56 14
rect -82 -68 -80 -48
rect -74 -68 -72 -48
rect -58 -68 -56 -48
rect -42 -68 -40 -48
rect -34 -68 -32 -48
rect 13 -67 15 -47
rect 21 -67 23 -47
rect 37 -67 39 -47
rect 53 -67 55 -47
rect 61 -67 63 -47
rect 77 -67 79 -47
<< ndiffusion >>
rect -67 -22 -66 -18
rect -71 -28 -66 -22
rect -64 -24 -58 -18
rect -64 -28 -63 -24
rect -59 -28 -58 -24
rect -56 -22 -55 -18
rect -56 -28 -51 -22
rect -83 -84 -82 -80
rect -87 -90 -82 -84
rect -80 -86 -74 -80
rect -80 -90 -79 -86
rect -75 -90 -74 -86
rect -72 -84 -71 -80
rect -72 -90 -67 -84
rect -63 -86 -58 -80
rect -59 -90 -58 -86
rect -56 -84 -55 -80
rect -56 -90 -51 -84
rect -47 -96 -42 -80
rect -43 -100 -42 -96
rect -40 -100 -34 -80
rect -32 -84 -31 -80
rect -32 -100 -27 -84
rect 8 -95 13 -79
rect 12 -99 13 -95
rect 15 -99 21 -79
rect 23 -83 24 -79
rect 23 -99 28 -83
rect 32 -85 37 -79
rect 36 -89 37 -85
rect 39 -83 40 -79
rect 39 -89 44 -83
rect 52 -83 53 -79
rect 48 -89 53 -83
rect 55 -85 61 -79
rect 55 -89 56 -85
rect 60 -89 61 -85
rect 63 -83 64 -79
rect 63 -89 68 -83
rect 72 -85 77 -79
rect 76 -89 77 -85
rect 79 -83 80 -79
rect 79 -89 84 -83
<< pdiffusion >>
rect -67 10 -66 14
rect -71 -6 -66 10
rect -64 -6 -58 14
rect -56 -2 -51 14
rect -56 -6 -55 -2
rect -83 -52 -82 -48
rect -87 -68 -82 -52
rect -80 -68 -74 -48
rect -72 -64 -67 -48
rect -72 -68 -71 -64
rect -59 -52 -58 -48
rect -63 -68 -58 -52
rect -56 -64 -51 -48
rect -56 -68 -55 -64
rect -43 -52 -42 -48
rect -47 -68 -42 -52
rect -40 -64 -34 -48
rect -40 -68 -39 -64
rect -35 -68 -34 -64
rect -32 -52 -31 -48
rect -32 -68 -27 -52
rect 12 -51 13 -47
rect 8 -67 13 -51
rect 15 -63 21 -47
rect 15 -67 16 -63
rect 20 -67 21 -63
rect 23 -51 24 -47
rect 23 -67 28 -51
rect 36 -51 37 -47
rect 32 -67 37 -51
rect 39 -63 44 -47
rect 39 -67 40 -63
rect 52 -51 53 -47
rect 48 -67 53 -51
rect 55 -67 61 -47
rect 63 -63 68 -47
rect 63 -67 64 -63
rect 76 -51 77 -47
rect 72 -67 77 -51
rect 79 -63 84 -47
rect 79 -67 80 -63
<< ndcontact >>
rect -71 -22 -67 -18
rect -63 -28 -59 -24
rect -55 -22 -51 -18
rect -87 -84 -83 -80
rect -79 -90 -75 -86
rect -71 -84 -67 -80
rect -63 -90 -59 -86
rect -55 -84 -51 -80
rect -47 -100 -43 -96
rect -31 -84 -27 -80
rect 8 -99 12 -95
rect 24 -83 28 -79
rect 32 -89 36 -85
rect 40 -83 44 -79
rect 48 -83 52 -79
rect 56 -89 60 -85
rect 64 -83 68 -79
rect 72 -89 76 -85
rect 80 -83 84 -79
<< pdcontact >>
rect -71 10 -67 14
rect -55 -6 -51 -2
rect -87 -52 -83 -48
rect -71 -68 -67 -64
rect -63 -52 -59 -48
rect -55 -68 -51 -64
rect -47 -52 -43 -48
rect -39 -68 -35 -64
rect -31 -52 -27 -48
rect 8 -51 12 -47
rect 16 -67 20 -63
rect 24 -51 28 -47
rect 32 -51 36 -47
rect 40 -67 44 -63
rect 48 -51 52 -47
rect 64 -67 68 -63
rect 72 -51 76 -47
rect 80 -67 84 -63
<< polysilicon >>
rect -66 14 -64 17
rect -58 14 -56 17
rect -66 -18 -64 -6
rect -58 -10 -56 -6
rect -58 -18 -56 -15
rect -66 -31 -64 -28
rect -58 -31 -56 -28
rect -82 -48 -80 -45
rect -74 -48 -72 -45
rect -58 -48 -56 -45
rect -42 -48 -40 -45
rect -34 -48 -32 -45
rect 13 -47 15 -44
rect 21 -47 23 -44
rect 37 -47 39 -44
rect 53 -47 55 -44
rect 61 -47 63 -44
rect 77 -47 79 -44
rect -82 -80 -80 -68
rect -74 -72 -72 -68
rect -74 -80 -72 -77
rect -58 -80 -56 -68
rect -42 -80 -40 -68
rect -34 -80 -32 -68
rect 13 -79 15 -67
rect 21 -79 23 -67
rect 37 -79 39 -67
rect 53 -79 55 -67
rect 61 -71 63 -67
rect 61 -79 63 -76
rect 77 -79 79 -67
rect -82 -93 -80 -90
rect -74 -93 -72 -90
rect -58 -93 -56 -90
rect 37 -92 39 -89
rect 53 -92 55 -89
rect 61 -92 63 -89
rect 77 -92 79 -89
rect -42 -103 -40 -100
rect -34 -102 -32 -100
rect 13 -102 15 -99
rect 21 -101 23 -99
<< polycontact >>
rect -70 -11 -66 -7
rect -86 -73 -82 -69
rect -62 -79 -58 -75
rect -46 -78 -42 -74
rect 9 -72 13 -68
rect 33 -72 37 -68
rect 49 -72 53 -68
rect 73 -78 77 -74
rect -36 -106 -32 -102
rect 19 -105 23 -101
<< metal1 >>
rect -77 18 -45 21
rect -71 14 -68 18
rect -51 -6 -47 -3
rect -78 -10 -70 -7
rect -50 -18 -47 -6
rect -67 -21 -55 -18
rect -51 -21 -47 -18
rect -62 -32 -59 -28
rect -71 -35 -50 -32
rect -93 -45 -21 -42
rect 2 -44 90 -41
rect -87 -48 -84 -45
rect -63 -48 -60 -45
rect -47 -48 -44 -45
rect -30 -48 -27 -45
rect 8 -47 11 -44
rect 25 -47 28 -44
rect 32 -47 35 -44
rect 48 -47 51 -44
rect 72 -47 75 -44
rect -67 -68 -63 -65
rect 68 -67 72 -64
rect -95 -72 -86 -69
rect -66 -75 -63 -68
rect -54 -75 -51 -68
rect -38 -70 -35 -68
rect -38 -73 -16 -70
rect -5 -72 9 -69
rect 17 -69 20 -67
rect 17 -72 33 -69
rect 41 -69 44 -67
rect 41 -72 49 -69
rect -66 -79 -62 -75
rect -54 -78 -46 -75
rect -66 -80 -63 -79
rect -54 -80 -51 -78
rect -83 -83 -71 -80
rect -67 -83 -63 -80
rect -27 -83 -24 -73
rect 25 -79 28 -72
rect 41 -79 44 -72
rect 69 -74 72 -67
rect 81 -74 84 -67
rect 69 -78 73 -74
rect 81 -77 96 -74
rect 69 -79 72 -78
rect 81 -79 84 -77
rect 52 -82 64 -79
rect 68 -82 72 -79
rect -78 -93 -75 -90
rect -63 -93 -60 -90
rect 32 -92 35 -89
rect 57 -92 60 -89
rect 72 -92 75 -89
rect -85 -96 -44 -93
rect 8 -95 75 -92
rect -95 -106 -36 -103
rect -4 -105 19 -102
<< pm12contact >>
rect -58 -15 -53 -10
rect -74 -77 -69 -72
rect 61 -76 66 -71
<< metal2 >>
rect -78 -15 -58 -12
rect -95 -77 -74 -74
rect -5 -76 61 -73
<< labels >>
rlabel metal1 14 -42 14 -42 5 VDD
rlabel metal1 41 -70 41 -70 3 A
rlabel metal1 52 -94 52 -94 1 gnd
rlabel metal1 54 -42 54 -42 5 VDD
rlabel metal1 82 -76 82 -76 1 out
rlabel metal1 -41 -43 -41 -43 5 VDD
rlabel metal1 -24 -72 -24 -72 1 out
rlabel metal1 -81 -43 -81 -43 5 VDD
rlabel metal1 -53 -77 -53 -77 1 out
rlabel metal1 -83 -95 -83 -95 1 gnd
rlabel metal1 -94 -105 -94 -105 3 interNAND
rlabel metal2 -94 -76 -94 -76 3 interORg
rlabel metal1 -94 -71 -94 -71 3 interORp
rlabel metal1 -4 -71 -4 -71 1 lastandC
rlabel metal1 -3 -104 -3 -104 1 lastandnr
rlabel metal2 -4 -75 -4 -75 1 lastORnd
rlabel metal1 -49 -14 -49 -14 7 out
rlabel metal2 -78 -14 -78 -14 3 B
rlabel metal1 -78 -9 -78 -9 3 A
rlabel metal1 -65 20 -65 20 5 VDD
rlabel metal1 -67 -34 -67 -34 1 gnd
<< end >>
