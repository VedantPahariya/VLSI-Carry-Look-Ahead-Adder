magic
tech scmos
timestamp 1731484135
<< nwell >>
rect -184 246 -152 283
rect -125 246 -101 259
rect -184 227 -101 246
rect -184 191 -125 227
rect -140 188 -125 191
rect -101 158 -81 199
<< ntransistor >>
rect -114 211 -112 221
rect -173 145 -171 185
rect -165 145 -163 185
rect -111 186 -107 188
rect -146 142 -144 182
rect -138 142 -136 182
rect -111 170 -107 172
<< ptransistor >>
rect -173 197 -171 277
rect -165 197 -163 277
rect -146 200 -144 240
rect -138 200 -136 240
rect -114 233 -112 253
rect -95 186 -87 188
rect -95 170 -87 172
<< ndiffusion >>
rect -119 215 -114 221
rect -115 211 -114 215
rect -112 217 -111 221
rect -112 211 -107 217
rect -174 181 -173 185
rect -178 145 -173 181
rect -171 149 -165 185
rect -171 145 -170 149
rect -166 145 -165 149
rect -163 181 -162 185
rect -111 188 -107 189
rect -111 185 -107 186
rect -163 145 -158 181
rect -151 146 -146 182
rect -147 142 -146 146
rect -144 142 -138 182
rect -136 178 -135 182
rect -136 142 -131 178
rect -111 172 -107 173
rect -111 169 -107 170
<< pdiffusion >>
rect -178 201 -173 277
rect -174 197 -173 201
rect -171 197 -165 277
rect -163 273 -162 277
rect -163 197 -158 273
rect -115 249 -114 253
rect -147 236 -146 240
rect -151 200 -146 236
rect -144 204 -138 240
rect -144 200 -143 204
rect -139 200 -138 204
rect -136 236 -135 240
rect -136 200 -131 236
rect -119 233 -114 249
rect -112 237 -107 253
rect -112 233 -111 237
rect -91 189 -87 193
rect -95 188 -87 189
rect -95 185 -87 186
rect -91 181 -87 185
rect -91 173 -87 177
rect -95 172 -87 173
rect -95 169 -87 170
rect -90 165 -87 169
<< ndcontact >>
rect -119 211 -115 215
rect -111 217 -107 221
rect -178 181 -174 185
rect -170 145 -166 149
rect -162 181 -158 185
rect -111 189 -107 193
rect -151 142 -147 146
rect -135 178 -131 182
rect -111 181 -107 185
rect -111 173 -107 177
<< pdcontact >>
rect -178 197 -174 201
rect -162 273 -158 277
rect -119 249 -115 253
rect -151 236 -147 240
rect -143 200 -139 204
rect -135 236 -131 240
rect -111 233 -107 237
rect -95 189 -91 193
rect -95 181 -91 185
rect -95 173 -91 177
<< polysilicon >>
rect -173 277 -171 280
rect -165 277 -163 280
rect -114 253 -112 256
rect -146 240 -144 243
rect -138 240 -136 243
rect -114 221 -112 233
rect -114 208 -112 211
rect -173 193 -171 197
rect -173 185 -171 188
rect -165 185 -163 197
rect -146 182 -144 200
rect -138 192 -136 200
rect -138 182 -136 187
rect -114 186 -111 188
rect -107 187 -104 188
rect -99 187 -95 188
rect -107 186 -95 187
rect -87 186 -84 188
rect -173 142 -171 145
rect -165 142 -163 145
rect -115 170 -111 172
rect -107 170 -104 172
rect -98 170 -95 172
rect -87 170 -86 172
rect -146 139 -144 142
rect -138 139 -136 142
<< polycontact >>
rect -118 222 -114 226
rect -163 192 -159 196
rect -150 192 -146 196
rect -119 170 -115 174
rect -86 170 -82 174
<< metal1 >>
rect -184 281 -151 284
rect -161 277 -158 281
rect -154 252 -151 281
rect -154 249 -119 252
rect -142 240 -139 249
rect -128 240 -91 243
rect -147 237 -135 240
rect -128 226 -125 240
rect -128 223 -118 226
rect -158 220 -125 223
rect -110 221 -107 233
rect -182 197 -178 200
rect -182 185 -179 197
rect -158 196 -155 220
rect -125 211 -119 214
rect -142 198 -139 200
rect -159 193 -150 196
rect -142 195 -128 198
rect -182 182 -178 185
rect -174 182 -162 185
rect -131 179 -128 195
rect -134 171 -131 178
rect -183 168 -131 171
rect -170 141 -167 145
rect -151 141 -147 142
rect -125 141 -122 211
rect -110 193 -107 217
rect -94 198 -91 240
rect -94 195 -83 198
rect -94 193 -91 195
rect -118 190 -111 193
rect -118 174 -115 190
rect -107 181 -95 184
rect -105 177 -102 181
rect -107 174 -95 177
rect -103 160 -100 174
rect -86 174 -83 195
rect -179 138 -122 141
<< pm12contact >>
rect -176 188 -171 193
rect -140 187 -135 192
rect -104 187 -99 192
<< pdm12contact >>
rect -95 164 -90 169
<< ndm12contact >>
rect -112 164 -107 169
<< metal2 >>
rect -171 188 -140 191
rect -135 188 -104 191
rect -102 168 -99 187
rect -107 165 -95 168
<< labels >>
rlabel metal2 -156 189 -156 189 7 B
rlabel metal1 -156 194 -156 194 7 A
rlabel metal1 -164 283 -164 283 5 VDD
rlabel metal1 -162 139 -162 139 1 gnd
rlabel metal1 -181 186 -181 186 3 outnor
rlabel metal1 -182 169 -182 169 3 outnand
rlabel metal1 -102 161 -102 161 1 outxor
<< end >>
