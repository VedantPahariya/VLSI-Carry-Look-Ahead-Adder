.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd

* Supply
Vdd vdd gnd 'SUPPLY'

* SPICE3 file created from TSPC3.ext - technology: scmos

.option scale=0.09u

M1000 gnd a_455_n375# a_451_n340# Gnd CMOSN w=20 l=2
+  ad=300 pd=160 as=80 ps=48
M1001 a_451_n340# clk Q Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1002 a_475_n340# clk a_455_n375# Gnd CMOSN w=20 l=2
+  ad=80 pd=48 as=100 ps=50
M1003 VDD a_479_n375# a_455_n375# w_444_n378# CMOSP w=20 l=2
+  ad=600 pd=280 as=100 ps=50
M1004 gnd D a_501_n395# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1005 gnd a_479_n375# a_475_n340# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 gnd a_501_n395# a_479_n375# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1007 a_497_n392# clk a_479_n375# w_444_n378# CMOSP w=40 l=2
+  ad=160 pd=88 as=200 ps=90
M1008 VDD D a_519_n392# w_444_n378# CMOSP w=40 l=2
+  ad=0 pd=0 as=160 ps=88
M1009 a_519_n392# clk a_501_n395# w_444_n378# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1010 VDD a_501_n395# a_497_n392# w_444_n378# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 VDD a_455_n375# Q w_444_n378# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
C0 Q a_519_n392# 0.01fF
C1 VDD a_519_n392# 0.01fF
C2 D a_501_n395# 0.05fF
C3 clk a_501_n395# 0.03fF
C4 clk a_479_n375# 0.33fF
C5 clk D 0.61fF
C6 Q a_497_n392# 0.01fF
C7 a_501_n395# w_444_n378# 0.09fF
C8 Q a_501_n395# 0.12fF
C9 w_444_n378# a_479_n375# 0.12fF
C10 D w_444_n378# 0.20fF
C11 Q a_479_n375# 0.12fF
C12 Q D 0.06fF
C13 VDD a_497_n392# 0.01fF
C14 gnd a_501_n395# 0.04fF
C15 gnd a_479_n375# 0.06fF
C16 gnd D 0.02fF
C17 clk w_444_n378# 0.37fF
C18 VDD a_501_n395# 0.08fF
C19 Q clk 0.19fF
C20 VDD a_479_n375# 0.08fF
C21 VDD D 0.06fF
C22 gnd a_451_n340# 0.01fF
C23 gnd clk 0.52fF
C24 Q w_444_n378# 0.14fF
C25 VDD clk 0.19fF
C26 gnd Q 0.02fF
C27 VDD w_444_n378# 0.12fF
C28 Q VDD 0.69fF
C29 clk a_455_n375# 0.09fF
C30 a_455_n375# w_444_n378# 0.11fF
C31 Q a_455_n375# 0.17fF
C32 gnd a_455_n375# 0.08fF
C33 gnd a_475_n340# 0.01fF
C34 VDD a_455_n375# 0.09fF
C35 VDD Gnd 0.03fF
C36 D Gnd 0.09fF
C37 a_501_n395# Gnd 0.15fF
C38 gnd Gnd 0.18fF
C39 Q Gnd 0.09fF
C40 a_479_n375# Gnd 0.10fF
C41 a_455_n375# Gnd 0.15fF
C42 clk Gnd 0.85fF
C43 w_444_n378# Gnd 4.00fF

V3 D gnd 'SUPPLY'
.ic V(Q) =0

.tran 0.1n 100n
V1 clk gnd PULSE 0 'SUPPLY' 30n 50p 50p 30n 60n
* V2 D gnd PULSE 0 'SUPPLY' 0 50p 50p 1.75n 3.5n

.control
run
plot V(Q) V(clk)+3 V(D)+6
.endc