.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd

* Supply
Vdd vdd gnd 'SUPPLY'

* SPICE3 file created from complete.ext - technology: scmos

.option scale=0.09u

M1000 gnd B_0 Pt0 Gnd CMOSN w=40 l=2
+  ad=4455 pd=2162 as=400 ps=180
M1001 a_44_n222# G0 gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1002 a_150_n274# C1 VDD w_137_n280# CMOSP w=20 l=2
+  ad=120 pd=52 as=8300 ps=3920
M1003 a_n101_n391# A_3 VDD w_n131_n463# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1004 a_174_n405# a_150_n383# VDD w_137_n389# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1005 a_190_n274# a_174_n296# VDD w_137_n280# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1006 S0 C0 pgxor0 w_38_n97# CMOSP w=8 l=2
+  ad=80 pd=52 as=120 ps=78
M1007 a_150_n165# C0 VDD w_137_n171# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1008 a_n30_n423# A_3 gnd Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1009 a_n101_n282# A_2 VDD w_n131_n354# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1010 a_190_n165# a_174_n187# VDD w_137_n171# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1011 C1 a_75_n113# VDD w_38_n97# CMOSP w=20 l=2
+  ad=160 pd=78 as=0 ps=0
M1012 a_44_n440# G2 a_51_n418# w_38_n424# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1013 a_n30_n314# A_2 gnd Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1014 a_174_n296# a_150_n274# VDD w_137_n280# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1015 a_195_n452# Pout gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1016 a_n101_n173# A_1 VDD w_n131_n245# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1017 gnd Pt3 P32 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1018 a_44_n222# G0 a_51_n200# w_38_n206# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1019 VDD G3 GPG3 w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1020 a_231_n296# C3 VDD w_137_n280# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1021 a_174_n187# a_150_n165# VDD w_137_n171# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1022 a_44_n331# G1 a_51_n309# w_38_n315# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1023 a_n30_n96# A_0 gnd Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1024 a_n30_n205# A_1 gnd Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1025 VDD G1 GPG1 w_38_n206# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1026 gnd a_174_n296# a_183_n296# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1027 gnd Pt2 P21 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1028 a_231_n187# C2 VDD w_137_n171# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1029 VDD G2 GPG2 w_38_n315# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1030 a_150_n383# P32 a_150_n415# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1031 gnd Pt1 P10 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1032 gnd a_174_n187# a_183_n187# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1033 a_44_n440# G2 gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1034 a_174_n296# a_150_n274# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1035 a_n101_n64# A_0 VDD w_n131_n136# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1036 a_150_n165# P10 a_150_n197# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1037 a_174_n405# a_150_n383# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1038 a_231_n296# C3 gnd Gnd CMOSN w=10 l=2
+  ad=70 pd=48 as=0 ps=0
M1039 a_150_n274# P21 a_150_n306# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1040 VDD B_0 G0 w_n131_n136# CMOSP w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1041 a_174_n187# a_150_n165# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1042 pgxor1 C1 S1 w_123_n108# CMOSP w=8 l=2
+  ad=125 pd=80 as=80 ps=52
M1043 a_231_n187# C2 gnd Gnd CMOSN w=10 l=2
+  ad=70 pd=48 as=0 ps=0
M1044 a_195_n452# Pout a_195_n460# w_189_n473# CMOSP w=40 l=2
+  ad=200 pd=90 as=240 ps=92
M1045 a_136_n124# C1 VDD w_123_n108# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1046 Gout GPG3 gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1047 a_51_n91# Pt0 VDD w_38_n97# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1048 pgxor0 B_0 a_n101_n64# Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=70 ps=48
M1049 VDD G0 C1 w_38_n97# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 pgxor1 a_136_n124# S1 Gnd CMOSN w=4 l=2
+  ad=69 pd=58 as=40 ps=36
M1051 VDD P32 a_150_n383# w_137_n389# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1052 a_91_n341# a_75_n331# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1053 C4 a_216_n386# a_257_n392# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1054 a_136_n124# C1 gnd Gnd CMOSN w=10 l=2
+  ad=70 pd=48 as=0 ps=0
M1055 a_91_n232# a_75_n222# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1056 pgxor0 B_0 A_0 w_n47_n53# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1057 VDD P21 a_150_n274# w_137_n280# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 gnd Pt0 a_44_n123# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1059 P32 Pt2 a_76_n374# w_38_n424# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1060 gnd C0bar a_195_n452# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1061 VDD a_216_n386# C4 w_137_n389# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1062 a_183_n296# GPG2 a_190_n274# w_137_n280# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1063 a_91_n123# a_75_n113# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1064 VDD P10 a_150_n165# w_137_n171# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 P21 Pt1 a_76_n265# w_38_n315# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1066 a_183_n187# GPG1 a_190_n165# w_137_n171# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1067 C3 a_183_n296# VDD w_137_n280# CMOSP w=20 l=2
+  ad=140 pd=76 as=0 ps=0
M1068 pgxor2 B_2 a_n101_n282# Gnd CMOSN w=4 l=2
+  ad=69 pd=58 as=70 ps=48
M1069 P10 Pt0 a_76_n156# w_38_n206# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1070 C2 a_183_n187# VDD w_137_n171# CMOSP w=20 l=2
+  ad=140 pd=76 as=0 ps=0
M1071 pgxor3 B_3 A_3 w_n47_n380# CMOSP w=8 l=2
+  ad=125 pd=80 as=40 ps=26
M1072 pgxor1 B_1 a_n101_n173# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=70 ps=48
M1073 Gout GPG3 a_198_n403# w_137_n389# CMOSP w=40 l=2
+  ad=200 pd=90 as=240 ps=92
M1074 a_183_n296# GPG2 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 a_44_n123# C0bar a_51_n91# w_38_n97# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1076 C0 a_84_n59# S0 Gnd CMOSN w=4 l=2
+  ad=29 pd=22 as=40 ps=36
M1077 pgxor2 a_231_n187# S2 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1078 G0 A_0 VDD w_n131_n136# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 a_183_n187# GPG1 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1080 pgxor2 B_2 A_2 w_n47_n271# CMOSP w=8 l=2
+  ad=125 pd=80 as=40 ps=26
M1081 a_216_n386# a_195_n452# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1082 pgxor3 C3 S3 w_137_n280# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=52
M1083 a_216_n386# a_195_n452# VDD w_189_n473# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1084 a_91_n450# a_75_n440# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1085 C3 a_183_n296# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1086 a_195_n460# C0bar VDD w_189_n473# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 VDD A_3 a_n125_n450# w_n131_n463# CMOSP w=80 l=2
+  ad=0 pd=0 as=480 ps=172
M1088 C0 pgxor0 S0 w_38_n97# CMOSP w=8 l=2
+  ad=45 pd=28 as=0 ps=0
M1089 pgxor1 B_1 A_1 w_n47_n162# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1090 pgxor2 C2 S2 w_137_n171# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=52
M1091 VDD B_3 G3 w_n131_n463# CMOSP w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1092 C0bar C0 VDD w_n131_n136# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1093 C2 a_183_n187# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1094 gnd a_174_n405# Gout Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 VDD A_2 a_n125_n341# w_n131_n354# CMOSP w=80 l=2
+  ad=0 pd=0 as=480 ps=172
M1096 S1 pgxor1 a_136_n124# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1097 VDD B_1 G1 w_n131_n245# CMOSP w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1098 Pt3 A_3 gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1099 VDD B_2 G2 w_n131_n354# CMOSP w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1100 VDD A_1 a_n125_n232# w_n131_n245# CMOSP w=80 l=2
+  ad=0 pd=0 as=480 ps=172
M1101 gnd Pt2 a_44_n331# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1102 gnd P10 a_156_n444# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1103 Pt2 A_2 gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1104 gnd Pt1 a_44_n222# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1105 a_257_n392# Gout gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 VDD A_0 a_n125_n123# w_n131_n136# CMOSP w=80 l=2
+  ad=0 pd=0 as=480 ps=172
M1107 pgxor3 B_3 a_n101_n391# Gnd CMOSN w=4 l=2
+  ad=69 pd=58 as=70 ps=48
M1108 C0bar C0 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1109 Pt1 A_1 gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1110 VDD P10 Pout w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1111 a_75_n331# a_44_n331# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1112 GPG2 G2 a_91_n341# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1113 a_76_n374# Pt3 VDD w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 Pt0 A_0 gnd Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 C4 Gout VDD w_137_n389# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 pgxor3 a_231_n296# S3 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1117 a_n101_n64# A_0 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1118 a_75_n222# a_44_n222# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1119 GPG1 G1 a_91_n232# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1120 a_51_n418# Pt3 VDD w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1121 a_44_n123# C0bar gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 a_76_n265# Pt2 VDD w_38_n315# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 B_2 a_n101_n282# pgxor2 Gnd CMOSN w=4 l=2
+  ad=29 pd=22 as=0 ps=0
M1124 a_51_n200# Pt1 VDD w_38_n206# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 G3 B_3 a_n30_n423# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1126 a_75_n113# a_44_n123# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1127 GPG3 a_75_n440# VDD w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 C1 G0 a_91_n123# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1129 a_76_n156# Pt1 VDD w_38_n206# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 a_51_n309# Pt2 VDD w_38_n315# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 G1 B_1 a_n30_n205# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1132 B_3 A_3 pgxor3 w_n47_n380# CMOSP w=8 l=2
+  ad=45 pd=28 as=0 ps=0
M1133 B_1 a_n101_n173# pgxor1 Gnd CMOSN w=4 l=2
+  ad=29 pd=22 as=0 ps=0
M1134 GPG1 a_75_n222# VDD w_38_n206# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 G2 B_2 a_n30_n314# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1136 S2 pgxor2 a_231_n187# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1137 a_75_n440# a_44_n440# VDD w_38_n424# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1138 GPG2 a_75_n331# VDD w_38_n315# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1139 a_198_n403# a_174_n405# VDD w_137_n389# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 P32 Pt2 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 S1 pgxor1 C1 w_123_n108# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 B_2 A_2 pgxor2 w_n47_n271# CMOSP w=8 l=2
+  ad=45 pd=28 as=0 ps=0
M1143 a_150_n415# GPG1 gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 G0 B_0 a_n30_n96# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1145 a_75_n222# a_44_n222# VDD w_38_n206# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1146 gnd Pt3 a_44_n440# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 S3 pgxor3 C3 w_137_n280# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 a_75_n331# a_44_n331# VDD w_38_n315# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1149 P21 Pt1 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 a_150_n197# C0 gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1151 a_150_n306# C1 gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1152 B_1 A_1 pgxor1 w_n47_n162# CMOSP w=8 l=2
+  ad=45 pd=28 as=0 ps=0
M1153 a_n125_n450# B_3 Pt3 w_n131_n463# CMOSP w=80 l=2
+  ad=0 pd=0 as=400 ps=170
M1154 S2 pgxor2 C2 w_137_n171# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 P10 Pt0 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1156 a_n101_n391# A_3 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1157 G3 A_3 VDD w_n131_n463# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 B_0 a_n101_n64# pgxor0 Gnd CMOSN w=4 l=2
+  ad=29 pd=22 as=0 ps=0
M1159 a_75_n440# a_44_n440# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1160 a_84_n59# pgxor0 VDD w_38_n97# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1161 GPG3 G3 a_91_n450# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1162 a_n125_n341# B_2 Pt2 w_n131_n354# CMOSP w=80 l=2
+  ad=0 pd=0 as=400 ps=170
M1163 gnd B_3 Pt3 Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 G2 A_2 VDD w_n131_n354# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 a_n101_n282# A_2 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 a_75_n113# a_44_n123# VDD w_38_n97# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1167 a_n125_n232# B_1 Pt1 w_n131_n245# CMOSP w=80 l=2
+  ad=0 pd=0 as=400 ps=170
M1168 a_156_n444# P32 Pout Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1169 gnd B_2 Pt2 Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 a_n101_n173# A_1 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 G1 A_1 VDD w_n131_n245# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 B_3 a_n101_n391# pgxor3 Gnd CMOSN w=4 l=2
+  ad=29 pd=22 as=0 ps=0
M1173 B_0 A_0 pgxor0 w_n47_n53# CMOSP w=8 l=2
+  ad=45 pd=28 as=0 ps=0
M1174 a_n125_n123# B_0 Pt0 w_n131_n136# CMOSP w=80 l=2
+  ad=0 pd=0 as=400 ps=170
M1175 a_44_n331# G1 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 a_84_n59# pgxor0 gnd Gnd CMOSN w=10 l=2
+  ad=70 pd=48 as=0 ps=0
M1177 gnd B_1 Pt1 Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 a_150_n383# GPG1 VDD w_137_n389# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 S0 C0 a_84_n59# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1180 Pout P32 VDD w_38_n424# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 S3 pgxor3 a_231_n296# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 gnd w_n131_n245# 0.03fF
C1 GPG1 P32 0.09fF
C2 S1 a_136_n124# 0.12fF
C3 gnd G0 1.58fF
C4 pgxor3 GPG1 0.05fF
C5 w_38_n315# a_44_n331# 0.10fF
C6 gnd Pt3 0.60fF
C7 B_1 G1 0.37fF
C8 Pt0 B_0 0.20fF
C9 pgxor2 G1 0.75fF
C10 gnd Pt2 0.43fF
C11 w_137_n280# P10 0.02fF
C12 VDD a_44_n440# 0.08fF
C13 C0bar a_195_n452# 0.10fF
C14 VDD Gout 0.12fF
C15 B_2 Pt2 0.20fF
C16 Pt1 P21 0.28fF
C17 C0 w_n131_n136# 0.13fF
C18 gnd a_n101_n64# 0.28fF
C19 A_1 a_n101_n173# 0.12fF
C20 gnd B_0 0.12fF
C21 w_137_n171# a_183_n187# 0.10fF
C22 gnd A_3 0.07fF
C23 G0 w_n131_n136# 0.06fF
C24 w_38_n315# P21 0.08fF
C25 w_137_n280# VDD 0.23fF
C26 G3 a_n30_n423# 0.02fF
C27 gnd a_75_n222# 0.06fF
C28 pgxor2 S2 0.50fF
C29 a_183_n296# C3 0.04fF
C30 C0bar a_n125_n232# 0.00fF
C31 Pt1 a_44_n222# 0.09fF
C32 w_n131_n245# B_1 0.44fF
C33 w_38_n206# P10 0.07fF
C34 G3 B_3 0.37fF
C35 a_n101_n64# w_n131_n136# 0.02fF
C36 w_n131_n354# G2 0.06fF
C37 A_2 Pt2 0.09fF
C38 pgxor1 C0 0.06fF
C39 a_183_n187# a_174_n187# 0.13fF
C40 B_0 w_n131_n136# 0.44fF
C41 C0bar a_n125_n123# 0.00fF
C42 gnd a_75_n113# 0.06fF
C43 VDD P10 0.19fF
C44 GPG1 a_150_n165# 0.07fF
C45 pgxor1 G0 0.75fF
C46 gnd a_183_n187# 0.12fF
C47 w_38_n206# VDD 0.16fF
C48 w_n131_n463# VDD 0.18fF
C49 pgxor3 w_137_n280# 0.37fF
C50 gnd a_n101_n173# 0.28fF
C51 a_75_n331# G2 0.09fF
C52 gnd a_195_n452# 0.18fF
C53 gnd G2 1.26fF
C54 P10 Pout 0.02fF
C55 w_n131_n463# a_n101_n391# 0.02fF
C56 B_2 G2 0.37fF
C57 gnd a_174_n296# 0.02fF
C58 a_44_n331# a_75_n331# 0.04fF
C59 a_174_n405# GPG3 0.14fF
C60 gnd a_44_n331# 0.12fF
C61 w_123_n108# C1 0.40fF
C62 a_150_n274# a_174_n296# 0.04fF
C63 P10 P32 0.46fF
C64 Pt3 w_38_n424# 0.25fF
C65 w_137_n171# GPG1 0.35fF
C66 VDD Pout 0.14fF
C67 GPG2 G2 0.06fF
C68 gnd G3 1.04fF
C69 pgxor3 P10 0.05fF
C70 gnd a_183_n296# 0.12fF
C71 gnd a_216_n386# 0.05fF
C72 Pt2 w_38_n424# 0.14fF
C73 w_137_n389# a_174_n405# 0.22fF
C74 GPG2 a_174_n296# 0.14fF
C75 w_38_n97# VDD 0.25fF
C76 C0 a_91_n123# 0.00fF
C77 C1 P21 0.09fF
C78 VDD P32 0.32fF
C79 a_44_n123# VDD 0.04fF
C80 gnd a_n125_n123# 0.01fF
C81 pgxor3 w_n47_n380# 0.07fF
C82 a_75_n440# G3 0.09fF
C83 G2 A_2 0.16fF
C84 pgxor3 VDD 0.24fF
C85 GPG1 C1 0.29fF
C86 C1 a_136_n124# 0.09fF
C87 gnd P21 0.29fF
C88 GPG1 a_174_n187# 0.14fF
C89 B_1 a_n101_n173# 0.20fF
C90 w_137_n389# C4 0.06fF
C91 GPG2 a_183_n296# 0.23fF
C92 C4 a_216_n386# 0.16fF
C93 Pt1 P10 0.14fF
C94 w_n131_n245# G1 0.06fF
C95 pgxor3 a_n101_n391# 0.12fF
C96 P21 a_150_n274# 0.06fF
C97 GPG1 gnd 0.18fF
C98 C2 VDD 0.09fF
C99 P32 Pout 0.15fF
C100 w_38_n206# Pt1 0.25fF
C101 pgxor1 a_n101_n173# 0.12fF
C102 w_137_n280# C3 0.27fF
C103 pgxor0 C0 0.29fF
C104 Pt2 G1 0.20fF
C105 GPG2 P21 0.17fF
C106 gnd a_44_n222# 0.12fF
C107 VDD Pt1 0.25fF
C108 a_44_n123# w_38_n97# 0.09fF
C109 w_n47_n53# C0bar 0.38fF
C110 GPG1 GPG2 0.05fF
C111 w_189_n473# a_195_n452# 0.10fF
C112 pgxor3 P32 0.46fF
C113 VDD w_38_n315# 0.16fF
C114 a_231_n296# S3 0.12fF
C115 a_150_n165# P10 0.06fF
C116 w_123_n108# pgxor1 0.41fF
C117 A_0 w_n47_n53# 0.19fF
C118 G1 a_75_n222# 0.09fF
C119 a_84_n59# pgxor0 0.23fF
C120 G0 C0 0.35fF
C121 gnd a_91_n232# 0.02fF
C122 G2 w_38_n424# 0.22fF
C123 pgxor0 a_n101_n64# 0.12fF
C124 pgxor2 P21 0.45fF
C125 pgxor0 B_0 0.52fF
C126 GPG3 w_38_n424# 0.30fF
C127 w_n131_n463# C0bar 0.20fF
C128 w_189_n473# a_216_n386# 0.03fF
C129 gnd a_44_n440# 0.12fF
C130 a_150_n165# VDD 0.02fF
C131 a_n101_n282# w_n131_n354# 0.02fF
C132 a_84_n59# C0 0.16fF
C133 GPG1 pgxor2 0.05fF
C134 gnd Gout 0.03fF
C135 w_n131_n463# B_3 0.44fF
C136 VDD C3 0.09fF
C137 Pt3 Pt2 0.07fF
C138 pgxor1 a_136_n124# 0.05fF
C139 VDD C0bar 1.23fF
C140 G3 w_38_n424# 0.06fF
C141 a_174_n405# Gout 0.09fF
C142 w_137_n280# C1 0.12fF
C143 w_n47_n380# B_3 0.28fF
C144 S0 pgxor0 0.10fF
C145 w_137_n171# P10 0.06fF
C146 w_n47_n162# A_1 0.19fF
C147 VDD B_3 0.06fF
C148 a_44_n440# a_75_n440# 0.04fF
C149 G0 B_0 0.37fF
C150 VDD A_1 0.28fF
C151 A_0 VDD 0.81fF
C152 a_n101_n282# gnd 0.28fF
C153 Pt3 A_3 0.09fF
C154 a_n101_n391# B_3 0.20fF
C155 GPG3 a_150_n383# 0.07fF
C156 C0bar Pout 0.08fF
C157 w_137_n280# a_150_n274# 0.15fF
C158 Gout C4 0.02fF
C159 a_n101_n282# B_2 0.20fF
C160 Pt0 P10 0.28fF
C161 S0 C0 0.50fF
C162 w_137_n171# VDD 0.23fF
C163 w_38_n206# Pt0 0.14fF
C164 w_137_n389# a_150_n383# 0.15fF
C165 w_38_n97# C0bar 0.21fF
C166 C1 P10 0.08fF
C167 C2 a_231_n187# 0.23fF
C168 w_137_n280# GPG2 0.35fF
C169 w_38_n315# Pt1 0.14fF
C170 a_44_n331# G1 0.06fF
C171 a_n101_n64# B_0 0.20fF
C172 VDD w_n131_n354# 0.18fF
C173 a_44_n123# C0bar 0.06fF
C174 pgxor3 C3 0.22fF
C175 C0 a_75_n113# 0.00fF
C176 gnd P10 0.47fF
C177 Pt0 VDD 0.21fF
C178 G0 a_75_n113# 0.09fF
C179 S0 a_84_n59# 0.12fF
C180 gnd w_n131_n463# 0.03fF
C181 pgxor3 B_3 0.52fF
C182 C1 VDD 0.22fF
C183 VDD a_174_n187# 0.02fF
C184 w_n131_n245# a_n101_n173# 0.02fF
C185 VDD a_75_n331# 0.08fF
C186 a_n101_n282# A_2 0.12fF
C187 gnd VDD 1.39fF
C188 GPG1 a_150_n383# 0.04fF
C189 GPG2 P10 0.05fF
C190 Pt3 G2 0.20fF
C191 VDD B_2 0.06fF
C192 VDD a_174_n405# 0.02fF
C193 VDD a_150_n274# 0.02fF
C194 Pt1 C0bar 0.00fF
C195 gnd a_n101_n391# 0.28fF
C196 a_n101_n282# pgxor2 0.12fF
C197 GPG1 G1 0.06fF
C198 Pt0 w_38_n97# 0.12fF
C199 G2 Pt2 0.85fF
C200 gnd Pout 0.19fF
C201 C2 w_137_n171# 0.27fF
C202 a_44_n123# Pt0 0.09fF
C203 VDD a_75_n440# 0.08fF
C204 Pt1 A_1 0.09fF
C205 gnd a_150_n306# 0.02fF
C206 gnd a_150_n415# 0.02fF
C207 C1 w_38_n97# 0.05fF
C208 VDD GPG2 0.04fF
C209 VDD C4 0.01fF
C210 C1 S1 0.11fF
C211 a_44_n440# w_38_n424# 0.10fF
C212 Pt3 G3 0.77fF
C213 VDD w_n131_n136# 0.24fF
C214 a_44_n331# Pt2 0.09fF
C215 gnd P32 0.32fF
C216 pgxor2 P10 0.08fF
C217 w_n47_n271# B_2 0.28fF
C218 a_44_n123# gnd 0.11fF
C219 pgxor3 gnd 0.90fF
C220 VDD A_2 0.28fF
C221 pgxor1 P10 0.29fF
C222 w_n47_n162# B_1 0.28fF
C223 GPG1 C0 0.04fF
C224 Pt0 Pt1 0.07fF
C225 VDD B_1 0.06fF
C226 C2 gnd 0.02fF
C227 G3 A_3 0.16fF
C228 pgxor2 VDD 0.24fF
C229 pgxor1 w_n47_n162# 0.07fF
C230 w_137_n171# a_231_n187# 0.02fF
C231 P21 Pt2 0.14fF
C232 C0bar B_3 0.00fF
C233 pgxor1 VDD 0.25fF
C234 C0bar A_1 0.00fF
C235 A_0 C0bar 0.10fF
C236 gnd Pt1 0.43fF
C237 w_137_n171# a_150_n165# 0.15fF
C238 G0 a_44_n222# 0.06fF
C239 w_n47_n271# A_2 0.19fF
C240 P10 w_38_n424# 0.17fF
C241 w_38_n315# a_75_n331# 0.10fF
C242 S3 w_137_n280# 0.06fF
C243 w_189_n473# VDD 0.07fF
C244 pgxor2 w_n47_n271# 0.07fF
C245 w_n131_n354# C0bar 0.20fF
C246 VDD w_38_n424# 0.26fF
C247 Pt0 C0bar 0.07fF
C248 a_150_n165# a_174_n187# 0.04fF
C249 w_189_n473# Pout 0.26fF
C250 pgxor1 S1 0.52fF
C251 w_38_n315# GPG2 0.19fF
C252 gnd a_150_n165# 0.04fF
C253 a_216_n386# a_195_n452# 0.04fF
C254 C2 pgxor2 0.22fF
C255 a_75_n222# a_44_n222# 0.04fF
C256 A_0 Pt0 0.09fF
C257 gnd C3 0.02fF
C258 gnd C0bar 0.47fF
C259 GPG3 G3 0.06fF
C260 w_38_n424# Pout 0.05fF
C261 pgxor0 w_n47_n53# 0.07fF
C262 Pt3 a_44_n440# 0.09fF
C263 w_137_n389# GPG3 0.50fF
C264 a_183_n296# a_174_n296# 0.13fF
C265 Pt1 B_1 0.20fF
C266 GPG1 a_183_n187# 0.23fF
C267 C0bar B_2 0.00fF
C268 w_38_n206# G1 0.06fF
C269 gnd B_3 0.11fF
C270 pgxor2 Pt1 0.27fF
C271 VDD a_150_n383# 0.02fF
C272 gnd A_1 0.07fF
C273 A_0 gnd 0.07fF
C274 w_137_n171# a_174_n187# 0.14fF
C275 w_137_n389# a_216_n386# 0.08fF
C276 w_38_n424# P32 0.19fF
C277 VDD G1 0.33fF
C278 C0bar w_n131_n136# 0.30fF
C279 GPG1 GPG3 0.00fF
C280 gnd w_n131_n354# 0.03fF
C281 pgxor2 a_231_n187# 0.16fF
C282 C0 P10 0.32fF
C283 pgxor0 VDD 0.46fF
C284 VDD a_51_n200# 0.01fF
C285 gnd Pt0 0.28fF
C286 A_0 w_n131_n136# 0.49fF
C287 w_n131_n354# B_2 0.44fF
C288 C0bar A_2 0.00fF
C289 GPG1 w_137_n389# 0.12fF
C290 P32 a_150_n383# 0.06fF
C291 w_123_n108# a_136_n124# 0.03fF
C292 gnd C1 0.27fF
C293 C0bar B_1 0.00fF
C294 gnd a_174_n187# 0.02fF
C295 w_38_n206# G0 0.22fF
C296 a_231_n296# w_137_n280# 0.02fF
C297 w_n47_n53# B_0 0.28fF
C298 gnd a_75_n331# 0.06fF
C299 pgxor3 S3 0.50fF
C300 w_n131_n463# Pt3 0.04fF
C301 C1 a_150_n274# 0.04fF
C302 VDD C0 3.15fF
C303 w_n131_n245# VDD 0.18fF
C304 A_1 B_1 0.32fF
C305 gnd B_2 0.11fF
C306 G0 VDD 0.29fF
C307 gnd a_174_n405# 0.06fF
C308 gnd a_150_n274# 0.04fF
C309 GPG1 P21 0.04fF
C310 VDD Pt3 0.14fF
C311 pgxor0 w_38_n97# 0.31fF
C312 Pt0 w_n131_n136# 0.04fF
C313 C1 GPG2 0.02fF
C314 a_44_n440# G2 0.06fF
C315 pgxor1 A_1 0.11fF
C316 VDD Pt2 0.25fF
C317 gnd a_150_n197# 0.02fF
C318 w_n131_n354# A_2 0.48fF
C319 w_137_n171# pgxor2 0.37fF
C320 VDD a_51_n309# 0.01fF
C321 w_189_n473# C0bar 0.18fF
C322 VDD a_51_n418# 0.01fF
C323 gnd GPG2 0.04fF
C324 a_84_n59# VDD 0.20fF
C325 w_n131_n463# A_3 0.48fF
C326 a_n30_n205# G1 0.02fF
C327 w_38_n206# a_75_n222# 0.10fF
C328 gnd w_n131_n136# 0.14fF
C329 a_51_n91# VDD 0.01fF
C330 w_38_n97# C0 0.95fF
C331 Pt1 G1 0.85fF
C332 GPG3 Gout 0.22fF
C333 VDD a_n101_n64# 0.02fF
C334 GPG2 a_150_n274# 0.07fF
C335 gnd a_91_n341# 0.02fF
C336 w_n47_n380# A_3 0.19fF
C337 VDD B_0 0.06fF
C338 a_44_n123# C0 0.07fF
C339 VDD A_3 0.28fF
C340 G0 w_38_n97# 0.06fF
C341 gnd a_156_n444# 0.02fF
C342 w_38_n315# G1 0.22fF
C343 VDD a_75_n222# 0.08fF
C344 gnd A_2 0.07fF
C345 C2 S2 0.10fF
C346 w_137_n389# Gout 0.23fF
C347 Pt3 P32 0.14fF
C348 a_n101_n391# A_3 0.12fF
C349 Pt0 pgxor1 0.27fF
C350 w_137_n280# a_174_n296# 0.14fF
C351 Gout a_216_n386# 0.31fF
C352 pgxor2 C1 0.36fF
C353 a_n125_n341# C0bar 0.00fF
C354 B_2 A_2 0.32fF
C355 gnd B_1 0.11fF
C356 Pt2 P32 0.28fF
C357 a_84_n59# w_38_n97# 0.02fF
C358 pgxor1 C1 0.77fF
C359 pgxor2 gnd 1.03fF
C360 pgxor3 Pt2 0.27fF
C361 w_137_n280# a_183_n296# 0.10fF
C362 pgxor2 B_2 0.52fF
C363 gnd pgxor1 0.96fF
C364 VDD a_195_n460# 0.02fF
C365 S3 C3 0.10fF
C366 VDD a_75_n113# 0.02fF
C367 w_n131_n245# Pt1 0.04fF
C368 a_183_n187# VDD 0.03fF
C369 GPG3 P10 0.05fF
C370 G0 Pt1 0.20fF
C371 pgxor3 A_3 0.11fF
C372 gnd w_189_n473# 0.10fF
C373 w_137_n280# P21 0.06fF
C374 Pout a_195_n460# 0.04fF
C375 VDD a_195_n452# 0.02fF
C376 a_231_n296# pgxor3 0.16fF
C377 S0 w_38_n97# 0.06fF
C378 VDD G2 0.33fF
C379 a_231_n187# S2 0.12fF
C380 a_n30_n96# G0 0.02fF
C381 Pt1 Pt2 0.07fF
C382 A_1 G1 0.16fF
C383 w_137_n389# P10 0.02fF
C384 pgxor0 C0bar 0.51fF
C385 VDD GPG3 0.07fF
C386 VDD a_174_n296# 0.02fF
C387 w_n131_n463# G3 0.06fF
C388 w_38_n315# Pt2 0.25fF
C389 w_38_n97# a_75_n113# 0.10fF
C390 pgxor2 A_2 0.11fF
C391 a_195_n452# Pout 0.22fF
C392 VDD a_44_n331# 0.08fF
C393 a_150_n165# C0 0.04fF
C394 a_44_n123# a_75_n113# 0.04fF
C395 A_0 pgxor0 0.11fF
C396 VDD G3 0.12fF
C397 w_137_n389# VDD 0.28fF
C398 w_123_n108# VDD 0.03fF
C399 P10 P21 0.04fF
C400 VDD a_183_n296# 0.03fF
C401 VDD a_216_n386# 0.06fF
C402 C0 C0bar 0.06fF
C403 pgxor1 B_1 0.52fF
C404 a_75_n440# w_38_n424# 0.10fF
C405 w_n131_n245# C0bar 0.20fF
C406 GPG1 P10 0.50fF
C407 G0 C0bar 0.02fF
C408 C2 a_183_n187# 0.04fF
C409 C0bar Pt3 0.00fF
C410 gnd a_150_n383# 0.04fF
C411 gnd a_91_n123# 0.02fF
C412 w_38_n206# GPG1 0.21fF
C413 pgxor3 G2 0.75fF
C414 w_n131_n245# A_1 0.48fF
C415 w_137_n171# S2 0.06fF
C416 GPG3 P32 0.17fF
C417 Pt3 B_3 0.20fF
C418 a_174_n405# a_150_n383# 0.04fF
C419 VDD P21 0.32fF
C420 C0bar Pt2 0.00fF
C421 A_0 G0 0.16fF
C422 gnd G1 1.26fF
C423 w_137_n171# C0 0.12fF
C424 C0bar a_n125_n450# 0.00fF
C425 GPG1 VDD 0.14fF
C426 w_38_n206# a_44_n222# 0.10fF
C427 w_137_n389# P32 0.06fF
C428 w_123_n108# S1 0.07fF
C429 B_0 C0bar 0.02fF
C430 C0bar A_3 0.00fF
C431 a_231_n296# C3 0.23fF
C432 gnd pgxor0 0.02fF
C433 Pt0 C0 0.01fF
C434 VDD a_44_n222# 0.08fF
C435 A_0 a_n101_n64# 0.12fF
C436 B_3 A_3 0.32fF
C437 A_0 B_0 0.32fF
C438 Pt0 G0 0.88fF
C439 C1 C0 0.11fF
C440 w_38_n315# G2 0.06fF
C441 w_n131_n354# Pt2 0.04fF
C442 G2 a_n30_n314# 0.02fF
C443 C1 G0 0.06fF
C444 gnd C0 0.30fF
C445 Pout Gnd 0.45fF
C446 a_195_n452# Gnd 0.16fF
C447 a_216_n386# Gnd 0.22fF
C448 C4 Gnd 0.06fF
C449 Gout Gnd 0.11fF
C450 G3 Gnd 0.43fF
C451 a_75_n440# Gnd 0.13fF
C452 a_44_n440# Gnd 0.02fF
C453 a_n101_n391# Gnd 0.26fF
C454 Pt3 Gnd 1.11fF
C455 GPG3 Gnd 0.92fF
C456 a_150_n383# Gnd 0.09fF
C457 P32 Gnd 0.60fF
C458 A_3 Gnd 0.43fF
C459 B_3 Gnd 0.74fF
C460 G2 Gnd 0.99fF
C461 a_75_n331# Gnd 0.13fF
C462 a_44_n331# Gnd 0.06fF
C463 a_n101_n282# Gnd 0.26fF
C464 S3 Gnd 0.08fF
C465 pgxor3 Gnd 2.60fF
C466 a_231_n296# Gnd 0.06fF
C467 Pt2 Gnd 1.65fF
C468 C3 Gnd 0.11fF
C469 a_183_n296# Gnd 0.15fF
C470 GPG2 Gnd 0.53fF
C471 a_174_n296# Gnd 0.09fF
C472 a_150_n274# Gnd 0.09fF
C473 P21 Gnd 0.05fF
C474 A_2 Gnd 0.43fF
C475 B_2 Gnd 0.74fF
C476 G1 Gnd 0.98fF
C477 a_75_n222# Gnd 0.13fF
C478 a_44_n222# Gnd 0.06fF
C479 a_n101_n173# Gnd 0.26fF
C480 S2 Gnd 0.08fF
C481 pgxor2 Gnd 2.56fF
C482 a_231_n187# Gnd 0.21fF
C483 Pt1 Gnd 1.65fF
C484 a_183_n187# Gnd 0.15fF
C485 GPG1 Gnd 1.38fF
C486 a_174_n187# Gnd 0.09fF
C487 a_150_n165# Gnd 0.09fF
C488 P10 Gnd 0.04fF
C489 A_1 Gnd 0.43fF
C490 B_1 Gnd 0.74fF
C491 S1 Gnd 0.12fF
C492 a_136_n124# Gnd 0.04fF
C493 pgxor1 Gnd 1.15fF
C494 C1 Gnd 0.55fF
C495 a_75_n113# Gnd 0.13fF
C496 G0 Gnd 0.00fF
C497 gnd Gnd 8.79fF
C498 a_n101_n64# Gnd 0.26fF
C499 Pt0 Gnd 1.37fF
C500 S0 Gnd 0.08fF
C501 a_84_n59# Gnd 0.21fF
C502 A_0 Gnd 0.42fF
C503 B_0 Gnd 0.74fF
C504 C0bar Gnd 8.27fF
C505 C0 Gnd 2.30fF
C506 VDD Gnd 0.01fF
C507 pgxor0 Gnd 0.43fF
C508 w_189_n473# Gnd 2.44fF
C509 w_137_n389# Gnd 4.21fF
C510 w_38_n424# Gnd 0.74fF
C511 w_n131_n463# Gnd 5.27fF
C512 w_n47_n380# Gnd 0.82fF
C513 w_137_n280# Gnd 0.01fF
C514 w_38_n315# Gnd 0.96fF
C515 w_n131_n354# Gnd 5.27fF
C516 w_n47_n271# Gnd 0.82fF
C517 w_137_n171# Gnd 0.39fF
C518 w_38_n206# Gnd 0.69fF
C519 w_n131_n245# Gnd 5.27fF
C520 w_n47_n162# Gnd 0.82fF
C521 w_123_n108# Gnd 0.31fF
C522 w_n47_n53# Gnd 0.82fF
C523 w_n131_n136# Gnd 6.10fF
C524 w_38_n97# Gnd 4.57fF


.tran 1n 10n

V1 A_0 gnd 'SUPPLY'
V2 A_1 gnd 0
V3 A_2 gnd 0
V4 A_3 gnd 0

V5 B_0 gnd 0
V6 B_1 gnd 0
V7 B_2 gnd 'SUPPLY'
V8 B_3 gnd 0
* V5 B_0 gnd PULSE(0 'SUPPLY' 50ns 50ps 50ps 30ns 60ns)
* V6 B1 gnd PULSE(0 'SUPPLY' 50ns 10ps 10ps 30ns 60ns)
* V7 B2 gnd PULSE(0 'SUPPLY' 50ns 10ps 10ps 30ns 60ns)

V9 C0 gnd 'SUPPLY'

.measure tran S0_val FIND v(S0) AT=8n
.measure tran S1_val FIND v(S1) AT=8n
.measure tran S2_val FIND v(S2) AT=8n  
.measure tran S3_val FIND v(S3) AT=8n  
.measure tran C4_val FIND v(C4) AT=8n
* .measure tran C1_val FIND v(C1) AT=8n
* .measure tran C2_val FIND v(C2) AT=8n
* .measure tran C3_val FIND v(C3) AT=8n
* .measure tran G0_val FIND v(G0) AT=8n
* .measure tran G2_val FIND v(G2) AT=8n
* .measure tran P2_val FIND v(Pt2) AT=8n
* .measure tran P21 FIND v(P21) AT=8n
* .measure tran P10 FIND v(P10) AT=8n
* .measure tran P1_val FIND v(Pt1) AT=8n
* .measure tran GPG2_val FIND v(GPG2) AT=8n
* .measure tran S2_val FIND v(S2) AT=16n
* .measure tran S3_val FIND v(S3) AT=16n
* .measure tran C4_val FIND v(Cout) AT=16n
 
.control
run
* plot V(S0)+3 V(S1) V(B_0)-3
.endc