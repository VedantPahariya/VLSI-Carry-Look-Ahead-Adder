magic
tech scmos
timestamp 1731446307
<< nwell >>
rect -209 29 -157 55
rect -42 40 -18 72
rect -7 42 25 74
rect 35 42 67 94
rect 76 42 108 134
rect -209 3 -108 29
rect -157 -3 -108 3
rect -123 -56 -78 -53
rect -143 -73 -78 -56
rect 21 -68 53 -13
rect 38 -71 53 -68
rect -143 -88 -119 -73
rect 96 -80 128 -45
rect 113 -83 128 -80
<< ntransistor >>
rect -145 35 -143 55
rect -139 35 -137 55
rect -121 35 -119 55
rect -115 35 -113 55
rect -31 24 -29 34
rect 4 26 6 36
rect 12 26 14 36
rect 46 16 48 36
rect 54 16 56 36
rect -198 -13 -196 -3
rect -176 -13 -174 -3
rect 87 -4 89 36
rect 95 -4 97 36
rect -108 -83 -106 -79
rect -92 -83 -90 -79
rect -132 -104 -130 -94
rect 32 -117 34 -77
rect 40 -117 42 -77
rect 107 -109 109 -89
rect 115 -109 117 -89
<< ptransistor >>
rect -198 9 -196 49
rect -192 9 -190 49
rect -176 9 -174 49
rect -170 9 -168 49
rect -31 46 -29 66
rect 4 48 6 68
rect 12 48 14 68
rect 46 48 48 88
rect 54 48 56 88
rect 87 48 89 128
rect 95 48 97 128
rect -145 3 -143 23
rect -121 3 -119 23
rect 32 -59 34 -19
rect 40 -59 42 -19
rect -132 -82 -130 -62
rect -108 -67 -106 -59
rect -92 -67 -90 -59
rect 107 -71 109 -51
rect 115 -71 117 -51
<< ndiffusion >>
rect -151 42 -145 55
rect -146 37 -145 42
rect -151 35 -145 37
rect -143 35 -139 55
rect -137 39 -131 55
rect -137 35 -135 39
rect -127 42 -121 55
rect -122 37 -121 42
rect -127 35 -121 37
rect -119 35 -115 55
rect -113 39 -107 55
rect -113 35 -111 39
rect -36 28 -31 34
rect -32 24 -31 28
rect -29 30 -28 34
rect -29 24 -24 30
rect 3 32 4 36
rect -1 26 4 32
rect 6 30 12 36
rect 6 26 7 30
rect 11 26 12 30
rect 14 32 15 36
rect 14 26 19 32
rect 45 32 46 36
rect 41 16 46 32
rect 48 20 54 36
rect 48 16 49 20
rect 53 16 54 20
rect 56 32 57 36
rect 56 16 61 32
rect 86 32 87 36
rect -203 -9 -198 -3
rect -199 -13 -198 -9
rect -196 -7 -195 -3
rect -196 -13 -191 -7
rect -181 -9 -176 -3
rect -177 -13 -176 -9
rect -174 -7 -173 -3
rect 82 -4 87 32
rect 89 0 95 36
rect 89 -4 90 0
rect 94 -4 95 0
rect 97 32 98 36
rect 97 -4 102 32
rect -174 -13 -169 -7
rect -109 -83 -108 -79
rect -106 -83 -105 -79
rect -93 -83 -92 -79
rect -90 -83 -89 -79
rect -137 -100 -132 -94
rect -133 -104 -132 -100
rect -130 -98 -129 -94
rect -130 -104 -125 -98
rect 27 -113 32 -77
rect 31 -117 32 -113
rect 34 -117 40 -77
rect 42 -81 43 -77
rect 42 -117 47 -81
rect 102 -105 107 -89
rect 106 -109 107 -105
rect 109 -109 115 -89
rect 117 -93 118 -89
rect 117 -109 122 -93
<< pdiffusion >>
rect 86 124 87 128
rect 45 84 46 88
rect -32 62 -31 66
rect -199 45 -198 49
rect -203 9 -198 45
rect -196 9 -192 49
rect -190 13 -185 49
rect -190 9 -189 13
rect -177 45 -176 49
rect -181 9 -176 45
rect -174 9 -170 49
rect -168 13 -163 49
rect -36 46 -31 62
rect -29 50 -24 66
rect -29 46 -28 50
rect 3 64 4 68
rect -1 48 4 64
rect 6 48 12 68
rect 14 52 19 68
rect 14 48 15 52
rect 41 48 46 84
rect 48 48 54 88
rect 56 52 61 88
rect 56 48 57 52
rect 82 48 87 124
rect 89 48 95 128
rect 97 52 102 128
rect 97 48 98 52
rect -168 9 -167 13
rect -150 9 -145 23
rect -146 5 -145 9
rect -150 3 -145 5
rect -143 19 -142 23
rect -143 3 -138 19
rect -126 9 -121 23
rect -122 5 -121 9
rect -126 3 -121 5
rect -119 19 -118 23
rect -119 3 -114 19
rect 31 -23 32 -19
rect 27 -59 32 -23
rect 34 -55 40 -19
rect 34 -59 35 -55
rect 39 -59 40 -55
rect 42 -23 43 -19
rect 42 -59 47 -23
rect 106 -55 107 -51
rect -133 -66 -132 -62
rect -137 -82 -132 -66
rect -130 -78 -125 -62
rect -113 -63 -108 -59
rect -109 -67 -108 -63
rect -106 -63 -101 -59
rect -106 -67 -105 -63
rect -97 -63 -92 -59
rect -93 -67 -92 -63
rect -90 -62 -85 -59
rect -90 -67 -89 -62
rect -130 -82 -129 -78
rect 102 -71 107 -55
rect 109 -67 115 -51
rect 109 -71 110 -67
rect 114 -71 115 -67
rect 117 -55 118 -51
rect 117 -71 122 -55
<< ndcontact >>
rect -135 35 -131 39
rect -111 35 -107 39
rect -36 24 -32 28
rect -28 30 -24 34
rect -1 32 3 36
rect 7 26 11 30
rect 15 32 19 36
rect 41 32 45 36
rect 49 16 53 20
rect 57 32 61 36
rect 82 32 86 36
rect -203 -13 -199 -9
rect -195 -7 -191 -3
rect -181 -13 -177 -9
rect -173 -7 -169 -3
rect 90 -4 94 0
rect 98 32 102 36
rect -113 -83 -109 -79
rect -105 -83 -101 -79
rect -97 -83 -93 -79
rect -137 -104 -133 -100
rect -129 -98 -125 -94
rect 27 -117 31 -113
rect 43 -81 47 -77
rect 102 -109 106 -105
rect 118 -93 122 -89
<< pdcontact >>
rect 82 124 86 128
rect 41 84 45 88
rect -36 62 -32 66
rect -203 45 -199 49
rect -189 9 -185 13
rect -181 45 -177 49
rect -28 46 -24 50
rect -1 64 3 68
rect 15 48 19 52
rect 57 48 61 52
rect 98 48 102 52
rect -167 9 -163 13
rect -150 5 -146 9
rect -142 19 -138 23
rect -126 5 -122 9
rect -118 19 -114 23
rect 27 -23 31 -19
rect 35 -59 39 -55
rect 43 -23 47 -19
rect 102 -55 106 -51
rect -137 -66 -133 -62
rect -113 -67 -109 -63
rect -105 -67 -101 -63
rect -97 -67 -93 -63
rect -129 -82 -125 -78
rect 110 -71 114 -67
rect 118 -55 122 -51
<< polysilicon >>
rect 87 128 89 131
rect 95 128 97 131
rect 46 88 48 91
rect 54 88 56 91
rect -31 66 -29 69
rect 4 68 6 71
rect 12 68 14 71
rect -198 49 -196 52
rect -192 49 -190 60
rect -176 49 -174 52
rect -170 49 -168 56
rect -145 55 -143 59
rect -139 55 -137 56
rect -121 55 -119 59
rect -115 55 -113 56
rect -145 23 -143 35
rect -139 32 -137 35
rect -121 23 -119 35
rect -115 32 -113 35
rect -31 34 -29 46
rect 4 36 6 48
rect 12 44 14 48
rect 12 36 14 39
rect 46 36 48 48
rect 54 44 56 48
rect 54 36 56 39
rect 87 36 89 48
rect 95 44 97 48
rect 95 36 97 39
rect -198 -3 -196 9
rect -192 6 -190 9
rect -176 -3 -174 9
rect -170 6 -168 9
rect -31 21 -29 24
rect 4 23 6 26
rect 12 23 14 26
rect 46 13 48 16
rect 54 13 56 16
rect -145 0 -143 3
rect -121 0 -119 3
rect 87 -7 89 -4
rect 95 -7 97 -4
rect -198 -16 -196 -13
rect -176 -16 -174 -13
rect 32 -19 34 -16
rect 40 -19 42 -16
rect -108 -59 -106 -56
rect -92 -59 -90 -58
rect 107 -51 109 -48
rect 115 -51 117 -48
rect -132 -62 -130 -59
rect -108 -71 -106 -67
rect -92 -70 -90 -67
rect -107 -76 -106 -71
rect -108 -79 -106 -76
rect -92 -79 -90 -76
rect 32 -77 34 -59
rect 40 -67 42 -59
rect 40 -77 42 -72
rect -132 -94 -130 -82
rect -108 -86 -106 -83
rect -92 -87 -90 -83
rect -132 -107 -130 -104
rect 107 -89 109 -71
rect 115 -79 117 -71
rect 115 -89 117 -84
rect 107 -112 109 -109
rect 115 -112 117 -109
rect 32 -120 34 -117
rect 40 -120 42 -117
<< polycontact >>
rect -190 56 -186 60
rect -171 56 -167 60
rect -139 56 -135 60
rect -115 56 -111 60
rect -35 35 -31 39
rect -125 30 -121 34
rect 0 43 4 47
rect 42 43 46 47
rect 83 43 87 47
rect -202 -2 -198 2
rect -180 -2 -176 2
rect -149 -2 -145 2
rect -94 -58 -90 -54
rect 28 -67 32 -63
rect -136 -93 -132 -89
rect -94 -91 -90 -87
rect 103 -79 107 -75
<< metal1 >>
rect 76 132 108 135
rect 82 128 85 132
rect 35 92 67 95
rect 41 88 44 92
rect -42 72 -18 75
rect -7 72 25 75
rect -36 66 -33 72
rect -1 68 2 72
rect -186 57 -171 60
rect -167 57 -139 60
rect -135 57 -115 60
rect -202 50 -154 53
rect -202 49 -199 50
rect -181 49 -177 50
rect -188 2 -185 9
rect -166 2 -163 9
rect -157 9 -154 50
rect 19 48 23 51
rect 61 48 65 51
rect 102 48 106 51
rect -41 36 -35 39
rect -134 33 -131 35
rect -134 30 -125 33
rect -110 33 -107 35
rect -27 34 -24 46
rect -9 44 0 47
rect 20 36 23 48
rect 33 44 42 47
rect 62 36 65 48
rect 74 44 83 47
rect 103 36 106 48
rect -110 30 -101 33
rect 3 33 15 36
rect 19 33 23 36
rect 45 33 57 36
rect 61 33 65 36
rect 86 33 98 36
rect 102 33 106 36
rect -134 23 -131 30
rect -110 23 -107 30
rect -138 20 -131 23
rect -114 20 -107 23
rect -36 21 -33 24
rect 8 22 11 26
rect -36 18 -24 21
rect -1 19 20 22
rect 50 12 53 16
rect 41 9 62 12
rect -157 6 -150 9
rect -146 6 -126 9
rect -208 -1 -202 2
rect -188 -1 -180 2
rect -188 -3 -185 -1
rect -166 -1 -149 2
rect -166 -3 -163 -1
rect -191 -6 -185 -3
rect -169 -6 -163 -3
rect 91 -8 94 -4
rect 82 -11 103 -8
rect -203 -16 -200 -13
rect -181 -16 -178 -13
rect 21 -15 53 -12
rect -203 -19 -169 -16
rect 27 -19 30 -15
rect 44 -19 47 -15
rect 96 -47 128 -44
rect 102 -51 105 -47
rect 119 -51 122 -47
rect -143 -56 -123 -53
rect -137 -62 -134 -56
rect -118 -58 -94 -55
rect -118 -63 -115 -58
rect 36 -61 39 -59
rect -118 -67 -113 -63
rect -118 -69 -115 -67
rect -155 -76 -151 -73
rect -142 -72 -115 -69
rect -142 -89 -139 -72
rect -104 -74 -101 -67
rect 19 -66 28 -63
rect 36 -64 54 -61
rect -97 -72 -94 -67
rect -97 -74 -80 -72
rect -104 -75 -80 -74
rect -104 -77 -94 -75
rect -104 -79 -101 -77
rect -128 -87 -125 -82
rect -97 -79 -94 -77
rect -113 -87 -110 -83
rect 47 -80 50 -64
rect 111 -73 114 -71
rect 94 -78 103 -75
rect 111 -76 129 -73
rect -142 -92 -136 -89
rect -128 -90 -94 -87
rect -128 -94 -125 -90
rect 122 -92 125 -76
rect -137 -107 -134 -104
rect -137 -110 -125 -107
rect 102 -113 105 -109
rect 102 -116 121 -113
rect 27 -121 30 -117
rect 27 -124 46 -121
<< m2contact >>
rect -67 -9 -59 -3
rect -169 -20 -164 -15
rect -151 -76 -146 -71
<< pm12contact >>
rect 12 39 17 44
rect 54 39 59 44
rect 95 39 100 44
rect -67 11 -59 17
rect -112 -76 -107 -71
rect 38 -72 43 -67
rect 113 -84 118 -79
<< pdm12contact >>
rect -67 1 -59 7
rect -89 -67 -84 -62
<< ndm12contact >>
rect -151 37 -146 42
rect -127 37 -122 42
rect -89 -84 -84 -79
<< metal2 >>
rect -146 38 -127 42
rect -151 33 -148 37
rect -135 36 -131 38
rect -9 39 12 42
rect 33 39 54 42
rect 74 39 95 42
rect -160 30 -148 33
rect -160 -16 -157 30
rect -164 -19 -157 -16
rect -88 -71 -85 -67
rect 19 -71 38 -68
rect -146 -76 -112 -73
rect -107 -74 -85 -71
rect -88 -79 -85 -74
rect 94 -83 113 -80
<< labels >>
rlabel metal1 -201 51 -201 51 1 VDD
rlabel metal1 -181 58 -181 58 5 clk
rlabel pm12contact -63 14 -63 14 7 poly_m1_m2
rlabel pdm12contact -64 4 -64 4 7 pdiff_m1_m2
rlabel m2contact -64 -6 -64 -6 7 m2contact
rlabel metal1 -206 0 -206 0 3 D
rlabel metal1 -102 31 -102 31 1 Q
rlabel metal1 -187 -18 -187 -18 1 gnd
rlabel metal1 -34 74 -34 74 5 VDD
rlabel metal1 -31 19 -31 19 1 gnd
rlabel metal1 21 40 21 40 7 out
rlabel metal2 -8 40 -8 40 3 B
rlabel metal1 -8 45 -8 45 3 A
rlabel metal1 5 74 5 74 5 VDD
rlabel metal1 3 20 3 20 1 gnd
rlabel metal1 63 40 63 40 7 out
rlabel metal2 34 40 34 40 3 B
rlabel metal1 34 45 34 45 3 A
rlabel metal1 47 94 47 94 5 VDD
rlabel metal1 45 10 45 10 1 gnd
rlabel metal1 104 40 104 40 7 out
rlabel metal2 75 40 75 40 3 B
rlabel metal1 75 45 75 45 3 A
rlabel metal1 88 134 88 134 5 VDD
rlabel metal1 86 -10 86 -10 1 gnd
rlabel metal1 33 -13 33 -13 5 VDD
rlabel metal2 20 -70 20 -70 3 B
rlabel metal1 20 -65 20 -65 3 A
rlabel metal1 34 -123 34 -123 1 gnd
rlabel metal1 50 -63 50 -63 1 out
rlabel metal2 95 -82 95 -82 3 B
rlabel metal1 95 -77 95 -77 3 A
rlabel metal1 125 -75 125 -75 1 out
rlabel metal1 108 -45 108 -45 5 VDD
rlabel metal1 109 -115 109 -115 1 gnd
rlabel metal1 -135 -54 -135 -54 5 VDD
rlabel metal1 -132 -109 -132 -109 1 gnd
rlabel metal1 -154 -75 -154 -75 1 B
rlabel metal1 -140 -91 -140 -91 1 A
rlabel metal1 -81 -74 -81 -74 1 out
<< end >>
